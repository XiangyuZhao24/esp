`timescale 1ps / 1ps
module fft_Mul_64Sx64S_86S_4(
          in2,
          in1,
          out1,
          clk,
          clr
);
   input [63:0] in2;
   input [63:0] in1;
   output [85:0] out1;
   input clk;
   input clr;
wire clk, clr, mul_34_17_n_0, mul_34_17_n_1, mul_34_17_n_2, mul_34_17_n_3,
     mul_34_17_n_4, mul_34_17_n_5, mul_34_17_n_6, mul_34_17_n_7, mul_34_17_n_8,
     mul_34_17_n_9, mul_34_17_n_10, mul_34_17_n_11, mul_34_17_n_12,
     mul_34_17_n_13, mul_34_17_n_14, mul_34_17_n_15, mul_34_17_n_16,
     mul_34_17_n_17, mul_34_17_n_18, mul_34_17_n_19, mul_34_17_n_20,
     mul_34_17_n_21, mul_34_17_n_22, mul_34_17_n_23, mul_34_17_n_24,
     mul_34_17_n_25, mul_34_17_n_26, mul_34_17_n_27, mul_34_17_n_28,
     mul_34_17_n_29, mul_34_17_n_30, mul_34_17_n_31, mul_34_17_n_32,
     mul_34_17_n_33, mul_34_17_n_34, mul_34_17_n_35, mul_34_17_n_36,
     mul_34_17_n_37, mul_34_17_n_38, mul_34_17_n_39, mul_34_17_n_40,
     mul_34_17_n_41, mul_34_17_n_42, mul_34_17_n_43, mul_34_17_n_44,
     mul_34_17_n_45, mul_34_17_n_46, mul_34_17_n_47, mul_34_17_n_48,
     mul_34_17_n_49, mul_34_17_n_50, mul_34_17_n_51, mul_34_17_n_52,
     mul_34_17_n_53, mul_34_17_n_54, mul_34_17_n_55, mul_34_17_n_56,
     mul_34_17_n_57, mul_34_17_n_58, mul_34_17_n_59, mul_34_17_n_60,
     mul_34_17_n_61, mul_34_17_n_62, mul_34_17_n_63, mul_34_17_n_64,
     mul_34_17_n_65, mul_34_17_n_66, mul_34_17_n_67, mul_34_17_n_68,
     mul_34_17_n_69, mul_34_17_n_70, mul_34_17_n_71, mul_34_17_n_72,
     mul_34_17_n_73, mul_34_17_n_74, mul_34_17_n_75, mul_34_17_n_76,
     mul_34_17_n_77, mul_34_17_n_78, mul_34_17_n_79, mul_34_17_n_80,
     mul_34_17_n_81, mul_34_17_n_82, mul_34_17_n_83, mul_34_17_n_84,
     mul_34_17_n_85, mul_34_17_n_86, mul_34_17_n_87, mul_34_17_n_88,
     mul_34_17_n_89, mul_34_17_n_90, mul_34_17_n_91, mul_34_17_n_92,
     mul_34_17_n_93, mul_34_17_n_94, mul_34_17_n_95, mul_34_17_n_96,
     mul_34_17_n_97, mul_34_17_n_98, mul_34_17_n_99, mul_34_17_n_100,
     mul_34_17_n_101, mul_34_17_n_102, mul_34_17_n_103, mul_34_17_n_104,
     mul_34_17_n_105, mul_34_17_n_106, mul_34_17_n_107, mul_34_17_n_108,
     mul_34_17_n_109, mul_34_17_n_110, mul_34_17_n_111, mul_34_17_n_112,
     mul_34_17_n_113, mul_34_17_n_114, mul_34_17_n_115, mul_34_17_n_117,
     mul_34_17_n_118, mul_34_17_n_119, mul_34_17_n_120, mul_34_17_n_121,
     mul_34_17_n_122, mul_34_17_n_123, mul_34_17_n_124, mul_34_17_n_125,
     mul_34_17_n_126, mul_34_17_n_127, mul_34_17_n_128, mul_34_17_n_129,
     mul_34_17_n_130, mul_34_17_n_131, mul_34_17_n_132, mul_34_17_n_133,
     mul_34_17_n_134, mul_34_17_n_135, mul_34_17_n_136, mul_34_17_n_137,
     mul_34_17_n_138, mul_34_17_n_139, mul_34_17_n_140, mul_34_17_n_141,
     mul_34_17_n_142, mul_34_17_n_143, mul_34_17_n_144, mul_34_17_n_145,
     mul_34_17_n_146, mul_34_17_n_147, mul_34_17_n_148, mul_34_17_n_149,
     mul_34_17_n_150, mul_34_17_n_151, mul_34_17_n_152, mul_34_17_n_154,
     mul_34_17_n_155, mul_34_17_n_156, mul_34_17_n_157, mul_34_17_n_158,
     mul_34_17_n_159, mul_34_17_n_160, mul_34_17_n_161, mul_34_17_n_162,
     mul_34_17_n_163, mul_34_17_n_164, mul_34_17_n_165, mul_34_17_n_166,
     mul_34_17_n_167, mul_34_17_n_168, mul_34_17_n_169, mul_34_17_n_170,
     mul_34_17_n_171, mul_34_17_n_172, mul_34_17_n_173, mul_34_17_n_174,
     mul_34_17_n_175, mul_34_17_n_176, mul_34_17_n_177, mul_34_17_n_178,
     mul_34_17_n_179, mul_34_17_n_180, mul_34_17_n_181, mul_34_17_n_182,
     mul_34_17_n_183, mul_34_17_n_184, mul_34_17_n_185, mul_34_17_n_186,
     mul_34_17_n_187, mul_34_17_n_188, mul_34_17_n_189, mul_34_17_n_190,
     mul_34_17_n_191, mul_34_17_n_192, mul_34_17_n_193, mul_34_17_n_194,
     mul_34_17_n_195, mul_34_17_n_196, mul_34_17_n_197, mul_34_17_n_198,
     mul_34_17_n_199, mul_34_17_n_200, mul_34_17_n_201, mul_34_17_n_202,
     mul_34_17_n_203, mul_34_17_n_204, mul_34_17_n_205, mul_34_17_n_206,
     mul_34_17_n_207, mul_34_17_n_209, mul_34_17_n_210, mul_34_17_n_211,
     mul_34_17_n_213, mul_34_17_n_215, mul_34_17_n_218, mul_34_17_n_219,
     mul_34_17_n_221, mul_34_17_n_223, mul_34_17_n_224, mul_34_17_n_225,
     mul_34_17_n_226, mul_34_17_n_227, mul_34_17_n_228, mul_34_17_n_229,
     mul_34_17_n_230, mul_34_17_n_231, mul_34_17_n_232, mul_34_17_n_233,
     mul_34_17_n_234, mul_34_17_n_235, mul_34_17_n_236, mul_34_17_n_237,
     mul_34_17_n_238, mul_34_17_n_239, mul_34_17_n_240, mul_34_17_n_241,
     mul_34_17_n_242, mul_34_17_n_243, mul_34_17_n_244, mul_34_17_n_246,
     mul_34_17_n_247, mul_34_17_n_249, mul_34_17_n_250, mul_34_17_n_251,
     mul_34_17_n_253, mul_34_17_n_254, mul_34_17_n_255, mul_34_17_n_256,
     mul_34_17_n_257, mul_34_17_n_259, mul_34_17_n_260, mul_34_17_n_261,
     mul_34_17_n_262, mul_34_17_n_263, mul_34_17_n_264, mul_34_17_n_265,
     mul_34_17_n_266, mul_34_17_n_267, mul_34_17_n_268, mul_34_17_n_269,
     mul_34_17_n_270, mul_34_17_n_271, mul_34_17_n_272, mul_34_17_n_273,
     mul_34_17_n_274, mul_34_17_n_275, mul_34_17_n_276, mul_34_17_n_277,
     mul_34_17_n_278, mul_34_17_n_279, mul_34_17_n_280, mul_34_17_n_281,
     mul_34_17_n_282, mul_34_17_n_283, mul_34_17_n_284, mul_34_17_n_285,
     mul_34_17_n_286, mul_34_17_n_287, mul_34_17_n_290, mul_34_17_n_291,
     mul_34_17_n_292, mul_34_17_n_294, mul_34_17_n_299, mul_34_17_n_300,
     mul_34_17_n_301, mul_34_17_n_302, mul_34_17_n_303, mul_34_17_n_304,
     mul_34_17_n_305, mul_34_17_n_306, mul_34_17_n_308, mul_34_17_n_309,
     mul_34_17_n_310, mul_34_17_n_311, mul_34_17_n_312, mul_34_17_n_313,
     mul_34_17_n_314, mul_34_17_n_315, mul_34_17_n_316, mul_34_17_n_317,
     mul_34_17_n_318, mul_34_17_n_319, mul_34_17_n_320, mul_34_17_n_321,
     mul_34_17_n_322, mul_34_17_n_323, mul_34_17_n_324, mul_34_17_n_325,
     mul_34_17_n_326, mul_34_17_n_327, mul_34_17_n_328, mul_34_17_n_329,
     mul_34_17_n_330, mul_34_17_n_331, mul_34_17_n_332, mul_34_17_n_333,
     mul_34_17_n_334, mul_34_17_n_335, mul_34_17_n_336, mul_34_17_n_337,
     mul_34_17_n_338, mul_34_17_n_339, mul_34_17_n_340, mul_34_17_n_341,
     mul_34_17_n_342, mul_34_17_n_343, mul_34_17_n_344, mul_34_17_n_345,
     mul_34_17_n_346, mul_34_17_n_347, mul_34_17_n_348, mul_34_17_n_349,
     mul_34_17_n_350, mul_34_17_n_351, mul_34_17_n_352, mul_34_17_n_353,
     mul_34_17_n_354, mul_34_17_n_355, mul_34_17_n_356, mul_34_17_n_357,
     mul_34_17_n_358, mul_34_17_n_359, mul_34_17_n_360, mul_34_17_n_361,
     mul_34_17_n_362, mul_34_17_n_363, mul_34_17_n_364, mul_34_17_n_365,
     mul_34_17_n_366, mul_34_17_n_367, mul_34_17_n_368, mul_34_17_n_369,
     mul_34_17_n_370, mul_34_17_n_371, mul_34_17_n_372, mul_34_17_n_373,
     mul_34_17_n_374, mul_34_17_n_375, mul_34_17_n_376, mul_34_17_n_377,
     mul_34_17_n_378, mul_34_17_n_379, mul_34_17_n_380, mul_34_17_n_381,
     mul_34_17_n_382, mul_34_17_n_383, mul_34_17_n_384, mul_34_17_n_385,
     mul_34_17_n_386, mul_34_17_n_387, mul_34_17_n_388, mul_34_17_n_389,
     mul_34_17_n_390, mul_34_17_n_391, mul_34_17_n_392, mul_34_17_n_393,
     mul_34_17_n_394, mul_34_17_n_395, mul_34_17_n_396, mul_34_17_n_397,
     mul_34_17_n_398, mul_34_17_n_399, mul_34_17_n_400, mul_34_17_n_401,
     mul_34_17_n_402, mul_34_17_n_403, mul_34_17_n_404, mul_34_17_n_405,
     mul_34_17_n_406, mul_34_17_n_407, mul_34_17_n_408, mul_34_17_n_409,
     mul_34_17_n_410, mul_34_17_n_411, mul_34_17_n_412, mul_34_17_n_413,
     mul_34_17_n_414, mul_34_17_n_415, mul_34_17_n_416, mul_34_17_n_417,
     mul_34_17_n_418, mul_34_17_n_419, mul_34_17_n_420, mul_34_17_n_421,
     mul_34_17_n_422, mul_34_17_n_423, mul_34_17_n_424, mul_34_17_n_425,
     mul_34_17_n_426, mul_34_17_n_427, mul_34_17_n_428, mul_34_17_n_429,
     mul_34_17_n_430, mul_34_17_n_431, mul_34_17_n_432, mul_34_17_n_433,
     mul_34_17_n_434, mul_34_17_n_435, mul_34_17_n_436, mul_34_17_n_437,
     mul_34_17_n_438, mul_34_17_n_439, mul_34_17_n_440, mul_34_17_n_441,
     mul_34_17_n_442, mul_34_17_n_443, mul_34_17_n_444, mul_34_17_n_445,
     mul_34_17_n_446, mul_34_17_n_447, mul_34_17_n_448, mul_34_17_n_449,
     mul_34_17_n_450, mul_34_17_n_451, mul_34_17_n_452, mul_34_17_n_453,
     mul_34_17_n_454, mul_34_17_n_455, mul_34_17_n_456, mul_34_17_n_457,
     mul_34_17_n_458, mul_34_17_n_459, mul_34_17_n_460, mul_34_17_n_461,
     mul_34_17_n_462, mul_34_17_n_463, mul_34_17_n_464, mul_34_17_n_465,
     mul_34_17_n_466, mul_34_17_n_467, mul_34_17_n_468, mul_34_17_n_469,
     mul_34_17_n_470, mul_34_17_n_471, mul_34_17_n_472, mul_34_17_n_473,
     mul_34_17_n_474, mul_34_17_n_475, mul_34_17_n_476, mul_34_17_n_477,
     mul_34_17_n_478, mul_34_17_n_479, mul_34_17_n_480, mul_34_17_n_481,
     mul_34_17_n_482, mul_34_17_n_483, mul_34_17_n_484, mul_34_17_n_485,
     mul_34_17_n_486, mul_34_17_n_487, mul_34_17_n_488, mul_34_17_n_489,
     mul_34_17_n_490, mul_34_17_n_491, mul_34_17_n_492, mul_34_17_n_493,
     mul_34_17_n_494, mul_34_17_n_495, mul_34_17_n_496, mul_34_17_n_497,
     mul_34_17_n_498, mul_34_17_n_499, mul_34_17_n_500, mul_34_17_n_501,
     mul_34_17_n_502, mul_34_17_n_503, mul_34_17_n_504, mul_34_17_n_505,
     mul_34_17_n_506, mul_34_17_n_507, mul_34_17_n_508, mul_34_17_n_509,
     mul_34_17_n_510, mul_34_17_n_511, mul_34_17_n_512, mul_34_17_n_513,
     mul_34_17_n_514, mul_34_17_n_515, mul_34_17_n_516, mul_34_17_n_517,
     mul_34_17_n_518, mul_34_17_n_519, mul_34_17_n_520, mul_34_17_n_521,
     mul_34_17_n_522, mul_34_17_n_523, mul_34_17_n_524, mul_34_17_n_525,
     mul_34_17_n_526, mul_34_17_n_527, mul_34_17_n_528, mul_34_17_n_529,
     mul_34_17_n_530, mul_34_17_n_531, mul_34_17_n_532, mul_34_17_n_533,
     mul_34_17_n_534, mul_34_17_n_535, mul_34_17_n_536, mul_34_17_n_537,
     mul_34_17_n_538, mul_34_17_n_539, mul_34_17_n_540, mul_34_17_n_541,
     mul_34_17_n_542, mul_34_17_n_543, mul_34_17_n_544, mul_34_17_n_545,
     mul_34_17_n_546, mul_34_17_n_547, mul_34_17_n_548, mul_34_17_n_549,
     mul_34_17_n_550, mul_34_17_n_551, mul_34_17_n_552, mul_34_17_n_553,
     mul_34_17_n_554, mul_34_17_n_555, mul_34_17_n_556, mul_34_17_n_557,
     mul_34_17_n_558, mul_34_17_n_559, mul_34_17_n_560, mul_34_17_n_561,
     mul_34_17_n_562, mul_34_17_n_563, mul_34_17_n_564, mul_34_17_n_565,
     mul_34_17_n_566, mul_34_17_n_567, mul_34_17_n_568, mul_34_17_n_569,
     mul_34_17_n_570, mul_34_17_n_571, mul_34_17_n_634, mul_34_17_n_635,
     mul_34_17_n_636, mul_34_17_n_637, mul_34_17_n_638, mul_34_17_n_639,
     mul_34_17_n_640, mul_34_17_n_641, mul_34_17_n_642, mul_34_17_n_643,
     mul_34_17_n_644, mul_34_17_n_645, mul_34_17_n_646, mul_34_17_n_647,
     mul_34_17_n_648, mul_34_17_n_649, mul_34_17_n_650, mul_34_17_n_651,
     mul_34_17_n_652, mul_34_17_n_653, mul_34_17_n_654, mul_34_17_n_655,
     mul_34_17_n_656, mul_34_17_n_657, mul_34_17_n_658, mul_34_17_n_659,
     mul_34_17_n_660, mul_34_17_n_661, mul_34_17_n_662, mul_34_17_n_663,
     mul_34_17_n_664, mul_34_17_n_665, mul_34_17_n_666, mul_34_17_n_667,
     mul_34_17_n_668, mul_34_17_n_669, mul_34_17_n_670, mul_34_17_n_671,
     mul_34_17_n_672, mul_34_17_n_673, mul_34_17_n_674, mul_34_17_n_675,
     mul_34_17_n_676, mul_34_17_n_677, mul_34_17_n_678, mul_34_17_n_679,
     mul_34_17_n_680, mul_34_17_n_681, mul_34_17_n_682, mul_34_17_n_683,
     mul_34_17_n_684, mul_34_17_n_685, mul_34_17_n_686, mul_34_17_n_687,
     mul_34_17_n_688, mul_34_17_n_689, mul_34_17_n_690, mul_34_17_n_691,
     mul_34_17_n_692, mul_34_17_n_693, mul_34_17_n_694, mul_34_17_n_695,
     mul_34_17_n_696, mul_34_17_n_697, mul_34_17_n_698, mul_34_17_n_699,
     mul_34_17_n_700, mul_34_17_n_701, mul_34_17_n_702, mul_34_17_n_703,
     mul_34_17_n_704, mul_34_17_n_705, mul_34_17_n_706, mul_34_17_n_707,
     mul_34_17_n_708, mul_34_17_n_709, mul_34_17_n_710, mul_34_17_n_711,
     mul_34_17_n_712, mul_34_17_n_713, mul_34_17_n_714, mul_34_17_n_715,
     mul_34_17_n_716, mul_34_17_n_717, mul_34_17_n_718, mul_34_17_n_719,
     mul_34_17_n_720, mul_34_17_n_721, mul_34_17_n_722, mul_34_17_n_723,
     mul_34_17_n_724, mul_34_17_n_725, mul_34_17_n_726, mul_34_17_n_727,
     mul_34_17_n_728, mul_34_17_n_729, mul_34_17_n_730, mul_34_17_n_731,
     mul_34_17_n_732, mul_34_17_n_733, mul_34_17_n_734, mul_34_17_n_735,
     mul_34_17_n_736, mul_34_17_n_737, mul_34_17_n_738, mul_34_17_n_739,
     mul_34_17_n_740, mul_34_17_n_741, mul_34_17_n_742, mul_34_17_n_743,
     mul_34_17_n_744, mul_34_17_n_745, mul_34_17_n_746, mul_34_17_n_747,
     mul_34_17_n_748, mul_34_17_n_749, mul_34_17_n_750, mul_34_17_n_751,
     mul_34_17_n_752, mul_34_17_n_753, mul_34_17_n_754, mul_34_17_n_755,
     mul_34_17_n_756, mul_34_17_n_757, mul_34_17_n_758, mul_34_17_n_759,
     mul_34_17_n_760, mul_34_17_n_761, mul_34_17_n_762, mul_34_17_n_763,
     mul_34_17_n_764, mul_34_17_n_765, mul_34_17_n_766, mul_34_17_n_767,
     mul_34_17_n_768, mul_34_17_n_769, mul_34_17_n_770, mul_34_17_n_771,
     mul_34_17_n_772, mul_34_17_n_773, mul_34_17_n_774, mul_34_17_n_775,
     mul_34_17_n_776, mul_34_17_n_777, mul_34_17_n_778, mul_34_17_n_779,
     mul_34_17_n_780, mul_34_17_n_781, mul_34_17_n_782, mul_34_17_n_783,
     mul_34_17_n_784, mul_34_17_n_785, mul_34_17_n_786, mul_34_17_n_787,
     mul_34_17_n_788, mul_34_17_n_789, mul_34_17_n_790, mul_34_17_n_791,
     mul_34_17_n_792, mul_34_17_n_793, mul_34_17_n_794, mul_34_17_n_795,
     mul_34_17_n_796, mul_34_17_n_797, mul_34_17_n_798, mul_34_17_n_799,
     mul_34_17_n_800, mul_34_17_n_801, mul_34_17_n_802, mul_34_17_n_803,
     mul_34_17_n_804, mul_34_17_n_805, mul_34_17_n_806, mul_34_17_n_807,
     mul_34_17_n_808, mul_34_17_n_809, mul_34_17_n_810, mul_34_17_n_811,
     mul_34_17_n_812, mul_34_17_n_813, mul_34_17_n_814, mul_34_17_n_815,
     mul_34_17_n_816, mul_34_17_n_817, mul_34_17_n_818, mul_34_17_n_819,
     mul_34_17_n_820, mul_34_17_n_821, mul_34_17_n_822, mul_34_17_n_823,
     mul_34_17_n_824, mul_34_17_n_825, mul_34_17_n_826, mul_34_17_n_827,
     mul_34_17_n_828, mul_34_17_n_829, mul_34_17_n_830, mul_34_17_n_831,
     mul_34_17_n_832, mul_34_17_n_833, mul_34_17_n_834, mul_34_17_n_835,
     mul_34_17_n_836, mul_34_17_n_837, mul_34_17_n_838, mul_34_17_n_839,
     mul_34_17_n_840, mul_34_17_n_841, mul_34_17_n_842, mul_34_17_n_843,
     mul_34_17_n_844, mul_34_17_n_845, mul_34_17_n_846, mul_34_17_n_847,
     mul_34_17_n_848, mul_34_17_n_849, mul_34_17_n_850, mul_34_17_n_851,
     mul_34_17_n_852, mul_34_17_n_853, mul_34_17_n_854, mul_34_17_n_855,
     mul_34_17_n_856, mul_34_17_n_857, mul_34_17_n_858, mul_34_17_n_859,
     mul_34_17_n_860, mul_34_17_n_861, mul_34_17_n_862, mul_34_17_n_863,
     mul_34_17_n_864, mul_34_17_n_865, mul_34_17_n_866, mul_34_17_n_867,
     mul_34_17_n_868, mul_34_17_n_869, mul_34_17_n_870, mul_34_17_n_871,
     mul_34_17_n_872, mul_34_17_n_873, mul_34_17_n_874, mul_34_17_n_875,
     mul_34_17_n_876, mul_34_17_n_877, mul_34_17_n_878, mul_34_17_n_879,
     mul_34_17_n_880, mul_34_17_n_881, mul_34_17_n_882, mul_34_17_n_883,
     mul_34_17_n_884, mul_34_17_n_885, mul_34_17_n_886, mul_34_17_n_887,
     mul_34_17_n_888, mul_34_17_n_889, mul_34_17_n_890, mul_34_17_n_891,
     mul_34_17_n_892, mul_34_17_n_893, mul_34_17_n_894, mul_34_17_n_895,
     mul_34_17_n_896, mul_34_17_n_897, mul_34_17_n_898, mul_34_17_n_899,
     mul_34_17_n_900, mul_34_17_n_901, mul_34_17_n_902, mul_34_17_n_903,
     mul_34_17_n_904, mul_34_17_n_905, mul_34_17_n_906, mul_34_17_n_907,
     mul_34_17_n_908, mul_34_17_n_909, mul_34_17_n_910, mul_34_17_n_911,
     mul_34_17_n_912, mul_34_17_n_913, mul_34_17_n_914, mul_34_17_n_915,
     mul_34_17_n_916, mul_34_17_n_917, mul_34_17_n_918, mul_34_17_n_919,
     mul_34_17_n_920, mul_34_17_n_921, mul_34_17_n_922, mul_34_17_n_923,
     mul_34_17_n_924, mul_34_17_n_925, mul_34_17_n_926, mul_34_17_n_927,
     mul_34_17_n_928, mul_34_17_n_929, mul_34_17_n_930, mul_34_17_n_931,
     mul_34_17_n_932, mul_34_17_n_933, mul_34_17_n_934, mul_34_17_n_935,
     mul_34_17_n_936, mul_34_17_n_937, mul_34_17_n_938, mul_34_17_n_939,
     mul_34_17_n_940, mul_34_17_n_941, mul_34_17_n_942, mul_34_17_n_943,
     mul_34_17_n_944, mul_34_17_n_945, mul_34_17_n_946, mul_34_17_n_947,
     mul_34_17_n_948, mul_34_17_n_949, mul_34_17_n_950, mul_34_17_n_951,
     mul_34_17_n_952, mul_34_17_n_953, mul_34_17_n_954, mul_34_17_n_955,
     mul_34_17_n_956, mul_34_17_n_957, mul_34_17_n_958, mul_34_17_n_959,
     mul_34_17_n_960, mul_34_17_n_961, mul_34_17_n_962, mul_34_17_n_963,
     mul_34_17_n_964, mul_34_17_n_965, mul_34_17_n_966, mul_34_17_n_967,
     mul_34_17_n_968, mul_34_17_n_969, mul_34_17_n_970, mul_34_17_n_971,
     mul_34_17_n_972, mul_34_17_n_973, mul_34_17_n_974, mul_34_17_n_975,
     mul_34_17_n_976, mul_34_17_n_977, mul_34_17_n_978, mul_34_17_n_979,
     mul_34_17_n_980, mul_34_17_n_981, mul_34_17_n_982, mul_34_17_n_983,
     mul_34_17_n_984, mul_34_17_n_985, mul_34_17_n_986, mul_34_17_n_987,
     mul_34_17_n_988, mul_34_17_n_989, mul_34_17_n_990, mul_34_17_n_991,
     mul_34_17_n_992, mul_34_17_n_993, mul_34_17_n_994, mul_34_17_n_995,
     mul_34_17_n_996, mul_34_17_n_997, mul_34_17_n_998, mul_34_17_n_999,
     mul_34_17_n_1000, mul_34_17_n_1001, mul_34_17_n_1002, mul_34_17_n_1003,
     mul_34_17_n_1004, mul_34_17_n_1005, mul_34_17_n_1006, mul_34_17_n_1007,
     mul_34_17_n_1008, mul_34_17_n_1009, mul_34_17_n_1010, mul_34_17_n_1011,
     mul_34_17_n_1012, mul_34_17_n_1013, mul_34_17_n_1014, mul_34_17_n_1015,
     mul_34_17_n_1016, mul_34_17_n_1017, mul_34_17_n_1018, mul_34_17_n_1019,
     mul_34_17_n_1020, mul_34_17_n_1021, mul_34_17_n_1022, mul_34_17_n_1023,
     mul_34_17_n_1024, mul_34_17_n_1025, mul_34_17_n_1026, mul_34_17_n_1027,
     mul_34_17_n_1028, mul_34_17_n_1029, mul_34_17_n_1030, mul_34_17_n_1031,
     mul_34_17_n_1032, mul_34_17_n_1033, mul_34_17_n_1034, mul_34_17_n_1035,
     mul_34_17_n_1036, mul_34_17_n_1037, mul_34_17_n_1038, mul_34_17_n_1039,
     mul_34_17_n_1040, mul_34_17_n_1041, mul_34_17_n_1042, mul_34_17_n_1043,
     mul_34_17_n_1044, mul_34_17_n_1045, mul_34_17_n_1046, mul_34_17_n_1047,
     mul_34_17_n_1048, mul_34_17_n_1049, mul_34_17_n_1050, mul_34_17_n_1051,
     mul_34_17_n_1052, mul_34_17_n_1053, mul_34_17_n_1054, mul_34_17_n_1055,
     mul_34_17_n_1056, mul_34_17_n_1057, mul_34_17_n_1058, mul_34_17_n_1059,
     mul_34_17_n_1060, mul_34_17_n_1061, mul_34_17_n_1062, mul_34_17_n_1063,
     mul_34_17_n_1064, mul_34_17_n_1065, mul_34_17_n_1066, mul_34_17_n_1067,
     mul_34_17_n_1068, mul_34_17_n_1069, mul_34_17_n_1070, mul_34_17_n_1071,
     mul_34_17_n_1072, mul_34_17_n_1073, mul_34_17_n_1074, mul_34_17_n_1075,
     mul_34_17_n_1076, mul_34_17_n_1077, mul_34_17_n_1078, mul_34_17_n_1079,
     mul_34_17_n_1080, mul_34_17_n_1081, mul_34_17_n_1082, mul_34_17_n_1083,
     mul_34_17_n_1084, mul_34_17_n_1085, mul_34_17_n_1086, mul_34_17_n_1087,
     mul_34_17_n_1088, mul_34_17_n_1089, mul_34_17_n_1090, mul_34_17_n_1091,
     mul_34_17_n_1092, mul_34_17_n_1093, mul_34_17_n_1094, mul_34_17_n_1095,
     mul_34_17_n_1096, mul_34_17_n_1097, mul_34_17_n_1098, mul_34_17_n_1099,
     mul_34_17_n_1100, mul_34_17_n_1101, mul_34_17_n_1102, mul_34_17_n_1103,
     mul_34_17_n_1104, mul_34_17_n_1105, mul_34_17_n_1106, mul_34_17_n_1107,
     mul_34_17_n_1108, mul_34_17_n_1109, mul_34_17_n_1110, mul_34_17_n_1111,
     mul_34_17_n_1112, mul_34_17_n_1113, mul_34_17_n_1114, mul_34_17_n_1115,
     mul_34_17_n_1116, mul_34_17_n_1117, mul_34_17_n_1118, mul_34_17_n_1119,
     mul_34_17_n_1120, mul_34_17_n_1121, mul_34_17_n_1122, mul_34_17_n_1123,
     mul_34_17_n_1124, mul_34_17_n_1125, mul_34_17_n_1126, mul_34_17_n_1127,
     mul_34_17_n_1128, mul_34_17_n_1129, mul_34_17_n_1130, mul_34_17_n_1131,
     mul_34_17_n_1132, mul_34_17_n_1133, mul_34_17_n_1134, mul_34_17_n_1135,
     mul_34_17_n_1136, mul_34_17_n_1137, mul_34_17_n_1138, mul_34_17_n_1139,
     mul_34_17_n_1140, mul_34_17_n_1141, mul_34_17_n_1142, mul_34_17_n_1143,
     mul_34_17_n_1144, mul_34_17_n_1145, mul_34_17_n_1146, mul_34_17_n_1147,
     mul_34_17_n_1148, mul_34_17_n_1149, mul_34_17_n_1150, mul_34_17_n_1151,
     mul_34_17_n_1152, mul_34_17_n_1153, mul_34_17_n_1154, mul_34_17_n_1155,
     mul_34_17_n_1156, mul_34_17_n_1157, mul_34_17_n_1158, mul_34_17_n_1159,
     mul_34_17_n_1160, mul_34_17_n_1161, mul_34_17_n_1162, mul_34_17_n_1163,
     mul_34_17_n_1164, mul_34_17_n_1165, mul_34_17_n_1166, mul_34_17_n_1167,
     mul_34_17_n_1168, mul_34_17_n_1169, mul_34_17_n_1170, mul_34_17_n_1171,
     mul_34_17_n_1172, mul_34_17_n_1173, mul_34_17_n_1174, mul_34_17_n_1175,
     mul_34_17_n_1176, mul_34_17_n_1177, mul_34_17_n_1178, mul_34_17_n_1179,
     mul_34_17_n_1180, mul_34_17_n_1181, mul_34_17_n_1182, mul_34_17_n_1183,
     mul_34_17_n_1184, mul_34_17_n_1185, mul_34_17_n_1186, mul_34_17_n_1187,
     mul_34_17_n_1188, mul_34_17_n_1189, mul_34_17_n_1190, mul_34_17_n_1191,
     mul_34_17_n_1192, mul_34_17_n_1193, mul_34_17_n_1194, mul_34_17_n_1195,
     mul_34_17_n_1196, mul_34_17_n_1197, mul_34_17_n_1198, mul_34_17_n_1199,
     mul_34_17_n_1200, mul_34_17_n_1201, mul_34_17_n_1202, mul_34_17_n_1203,
     mul_34_17_n_1204, mul_34_17_n_1205, mul_34_17_n_1206, mul_34_17_n_1207,
     mul_34_17_n_1208, mul_34_17_n_1209, mul_34_17_n_1210, mul_34_17_n_1211,
     mul_34_17_n_1212, mul_34_17_n_1213, mul_34_17_n_1214, mul_34_17_n_1215,
     mul_34_17_n_1216, mul_34_17_n_1217, mul_34_17_n_1218, mul_34_17_n_1219,
     mul_34_17_n_1220, mul_34_17_n_1221, mul_34_17_n_1222, mul_34_17_n_1223,
     mul_34_17_n_1224, mul_34_17_n_1225, mul_34_17_n_1226, mul_34_17_n_1227,
     mul_34_17_n_1228, mul_34_17_n_1229, mul_34_17_n_1230, mul_34_17_n_1231,
     mul_34_17_n_1232, mul_34_17_n_1233, mul_34_17_n_1234, mul_34_17_n_1235,
     mul_34_17_n_1236, mul_34_17_n_1237, mul_34_17_n_1238, mul_34_17_n_1239,
     mul_34_17_n_1240, mul_34_17_n_1241, mul_34_17_n_1242, mul_34_17_n_1243,
     mul_34_17_n_1244, mul_34_17_n_1245, mul_34_17_n_1246, mul_34_17_n_1247,
     mul_34_17_n_1248, mul_34_17_n_1249, mul_34_17_n_1250, mul_34_17_n_1251,
     mul_34_17_n_1252, mul_34_17_n_1253, mul_34_17_n_1254, mul_34_17_n_1255,
     mul_34_17_n_1256, mul_34_17_n_1257, mul_34_17_n_1258, mul_34_17_n_1259,
     mul_34_17_n_1260, mul_34_17_n_1261, mul_34_17_n_1262, mul_34_17_n_1263,
     mul_34_17_n_1264, mul_34_17_n_1265, mul_34_17_n_1266, mul_34_17_n_1267,
     mul_34_17_n_1268, mul_34_17_n_1269, mul_34_17_n_1270, mul_34_17_n_1271,
     mul_34_17_n_1272, mul_34_17_n_1273, mul_34_17_n_1274, mul_34_17_n_1275,
     mul_34_17_n_1276, mul_34_17_n_1277, mul_34_17_n_1278, mul_34_17_n_1279,
     mul_34_17_n_1280, mul_34_17_n_1281, mul_34_17_n_1282, mul_34_17_n_1283,
     mul_34_17_n_1284, mul_34_17_n_1285, mul_34_17_n_1286, mul_34_17_n_1287,
     mul_34_17_n_1288, mul_34_17_n_1289, mul_34_17_n_1290, mul_34_17_n_1291,
     mul_34_17_n_1292, mul_34_17_n_1293, mul_34_17_n_1294, mul_34_17_n_1295,
     mul_34_17_n_1296, mul_34_17_n_1297, mul_34_17_n_1298, mul_34_17_n_1299,
     mul_34_17_n_1300, mul_34_17_n_1301, mul_34_17_n_1302, mul_34_17_n_1303,
     mul_34_17_n_1304, mul_34_17_n_1305, mul_34_17_n_1306, mul_34_17_n_1307,
     mul_34_17_n_1308, mul_34_17_n_1309, mul_34_17_n_1310, mul_34_17_n_1311,
     mul_34_17_n_1312, mul_34_17_n_1313, mul_34_17_n_1314, mul_34_17_n_1315,
     mul_34_17_n_1316, mul_34_17_n_1317, mul_34_17_n_1318, mul_34_17_n_1319,
     mul_34_17_n_1320, mul_34_17_n_1321, mul_34_17_n_1322, mul_34_17_n_1323,
     mul_34_17_n_1324, mul_34_17_n_1325, mul_34_17_n_1326, mul_34_17_n_1327,
     mul_34_17_n_1328, mul_34_17_n_1329, mul_34_17_n_1330, mul_34_17_n_1331,
     mul_34_17_n_1332, mul_34_17_n_1333, mul_34_17_n_1334, mul_34_17_n_1335,
     mul_34_17_n_1336, mul_34_17_n_1337, mul_34_17_n_1338, mul_34_17_n_1339,
     mul_34_17_n_1340, mul_34_17_n_1341, mul_34_17_n_1342, mul_34_17_n_1343,
     mul_34_17_n_1344, mul_34_17_n_1345, mul_34_17_n_1346, mul_34_17_n_1347,
     mul_34_17_n_1348, mul_34_17_n_1349, mul_34_17_n_1350, mul_34_17_n_1351,
     mul_34_17_n_1352, mul_34_17_n_1353, mul_34_17_n_1354, mul_34_17_n_1355,
     mul_34_17_n_1356, mul_34_17_n_1357, mul_34_17_n_1358, mul_34_17_n_1359,
     mul_34_17_n_1360, mul_34_17_n_1361, mul_34_17_n_1362, mul_34_17_n_1363,
     mul_34_17_n_1364, mul_34_17_n_1365, mul_34_17_n_1366, mul_34_17_n_1367,
     mul_34_17_n_1368, mul_34_17_n_1369, mul_34_17_n_1370, mul_34_17_n_1371,
     mul_34_17_n_1372, mul_34_17_n_1373, mul_34_17_n_1374, mul_34_17_n_1375,
     mul_34_17_n_1376, mul_34_17_n_1377, mul_34_17_n_1378, mul_34_17_n_1379,
     mul_34_17_n_1380, mul_34_17_n_1381, mul_34_17_n_1382, mul_34_17_n_1383,
     mul_34_17_n_1384, mul_34_17_n_1385, mul_34_17_n_1386, mul_34_17_n_1387,
     mul_34_17_n_1388, mul_34_17_n_1389, mul_34_17_n_1390, mul_34_17_n_1391,
     mul_34_17_n_1392, mul_34_17_n_1393, mul_34_17_n_1394, mul_34_17_n_1395,
     mul_34_17_n_1396, mul_34_17_n_1397, mul_34_17_n_1398, mul_34_17_n_1399,
     mul_34_17_n_1400, mul_34_17_n_1401, mul_34_17_n_1402, mul_34_17_n_1403,
     mul_34_17_n_1404, mul_34_17_n_1405, mul_34_17_n_1406, mul_34_17_n_1407,
     mul_34_17_n_1408, mul_34_17_n_1409, mul_34_17_n_1410, mul_34_17_n_1411,
     mul_34_17_n_1412, mul_34_17_n_1413, mul_34_17_n_1414, mul_34_17_n_1415,
     mul_34_17_n_1416, mul_34_17_n_1417, mul_34_17_n_1418, mul_34_17_n_1419,
     mul_34_17_n_1420, mul_34_17_n_1421, mul_34_17_n_1422, mul_34_17_n_1423,
     mul_34_17_n_1424, mul_34_17_n_1425, mul_34_17_n_1426, mul_34_17_n_1427,
     mul_34_17_n_1428, mul_34_17_n_1429, mul_34_17_n_1430, mul_34_17_n_1431,
     mul_34_17_n_1432, mul_34_17_n_1433, mul_34_17_n_1434, mul_34_17_n_1435,
     mul_34_17_n_1436, mul_34_17_n_1437, mul_34_17_n_1438, mul_34_17_n_1439,
     mul_34_17_n_1440, mul_34_17_n_1441, mul_34_17_n_1442, mul_34_17_n_1443,
     mul_34_17_n_1444, mul_34_17_n_1445, mul_34_17_n_1446, mul_34_17_n_1447,
     mul_34_17_n_1448, mul_34_17_n_1449, mul_34_17_n_1450, mul_34_17_n_1451,
     mul_34_17_n_1452, mul_34_17_n_1453, mul_34_17_n_1454, mul_34_17_n_1455,
     mul_34_17_n_1456, mul_34_17_n_1457, mul_34_17_n_1458, mul_34_17_n_1459,
     mul_34_17_n_1460, mul_34_17_n_1461, mul_34_17_n_1462, mul_34_17_n_1463,
     mul_34_17_n_1464, mul_34_17_n_1465, mul_34_17_n_1466, mul_34_17_n_1467,
     mul_34_17_n_1468, mul_34_17_n_1469, mul_34_17_n_1470, mul_34_17_n_1471,
     mul_34_17_n_1472, mul_34_17_n_1473, mul_34_17_n_1474, mul_34_17_n_1475,
     mul_34_17_n_1476, mul_34_17_n_1477, mul_34_17_n_1478, mul_34_17_n_1479,
     mul_34_17_n_1480, mul_34_17_n_1481, mul_34_17_n_1482, mul_34_17_n_1483,
     mul_34_17_n_1484, mul_34_17_n_1485, mul_34_17_n_1486, mul_34_17_n_1487,
     mul_34_17_n_1488, mul_34_17_n_1489, mul_34_17_n_1490, mul_34_17_n_1491,
     mul_34_17_n_1492, mul_34_17_n_1493, mul_34_17_n_1494, mul_34_17_n_1495,
     mul_34_17_n_1496, mul_34_17_n_1497, mul_34_17_n_1498, mul_34_17_n_1499,
     mul_34_17_n_1500, mul_34_17_n_1501, mul_34_17_n_1502, mul_34_17_n_1503,
     mul_34_17_n_1504, mul_34_17_n_1505, mul_34_17_n_1506, mul_34_17_n_1507,
     mul_34_17_n_1508, mul_34_17_n_1509, mul_34_17_n_1510, mul_34_17_n_1511,
     mul_34_17_n_1512, mul_34_17_n_1513, mul_34_17_n_1514, mul_34_17_n_1515,
     mul_34_17_n_1516, mul_34_17_n_1517, mul_34_17_n_1518, mul_34_17_n_1519,
     mul_34_17_n_1520, mul_34_17_n_1521, mul_34_17_n_1522, mul_34_17_n_1523,
     mul_34_17_n_1524, mul_34_17_n_1525, mul_34_17_n_1526, mul_34_17_n_1527,
     mul_34_17_n_1528, mul_34_17_n_1529, mul_34_17_n_1530, mul_34_17_n_1531,
     mul_34_17_n_1532, mul_34_17_n_1533, mul_34_17_n_1534, mul_34_17_n_1535,
     mul_34_17_n_1536, mul_34_17_n_1537, mul_34_17_n_1538, mul_34_17_n_1539,
     mul_34_17_n_1540, mul_34_17_n_1541, mul_34_17_n_1542, mul_34_17_n_1543,
     mul_34_17_n_1544, mul_34_17_n_1545, mul_34_17_n_1546, mul_34_17_n_1547,
     mul_34_17_n_1548, mul_34_17_n_1549, mul_34_17_n_1550, mul_34_17_n_1551,
     mul_34_17_n_1552, mul_34_17_n_1553, mul_34_17_n_1554, mul_34_17_n_1555,
     mul_34_17_n_1556, mul_34_17_n_1557, mul_34_17_n_1558, mul_34_17_n_1559,
     mul_34_17_n_1560, mul_34_17_n_1561, mul_34_17_n_1562, mul_34_17_n_1563,
     mul_34_17_n_1564, mul_34_17_n_1565, mul_34_17_n_1566, mul_34_17_n_1567,
     mul_34_17_n_1568, mul_34_17_n_1569, mul_34_17_n_1570, mul_34_17_n_1571,
     mul_34_17_n_1572, mul_34_17_n_1573, mul_34_17_n_1574, mul_34_17_n_1575,
     mul_34_17_n_1576, mul_34_17_n_1577, mul_34_17_n_1578, mul_34_17_n_1579,
     mul_34_17_n_1580, mul_34_17_n_1581, mul_34_17_n_1582, mul_34_17_n_1583,
     mul_34_17_n_1584, mul_34_17_n_1585, mul_34_17_n_1586, mul_34_17_n_1587,
     mul_34_17_n_1588, mul_34_17_n_1589, mul_34_17_n_1590, mul_34_17_n_1591,
     mul_34_17_n_1592, mul_34_17_n_1593, mul_34_17_n_1594, mul_34_17_n_1595,
     mul_34_17_n_1596, mul_34_17_n_1597, mul_34_17_n_1598, mul_34_17_n_1599,
     mul_34_17_n_1600, mul_34_17_n_1601, mul_34_17_n_1602, mul_34_17_n_1603,
     mul_34_17_n_1604, mul_34_17_n_1605, mul_34_17_n_1606, mul_34_17_n_1607,
     mul_34_17_n_1608, mul_34_17_n_1609, mul_34_17_n_1610, mul_34_17_n_1611,
     mul_34_17_n_1612, mul_34_17_n_1613, mul_34_17_n_1614, mul_34_17_n_1615,
     mul_34_17_n_1616, mul_34_17_n_1617, mul_34_17_n_1618, mul_34_17_n_1619,
     mul_34_17_n_1620, mul_34_17_n_1621, mul_34_17_n_1622, mul_34_17_n_1623,
     mul_34_17_n_1624, mul_34_17_n_1625, mul_34_17_n_1626, mul_34_17_n_1627,
     mul_34_17_n_1628, mul_34_17_n_1629, mul_34_17_n_1630, mul_34_17_n_1631,
     mul_34_17_n_1632, mul_34_17_n_1633, mul_34_17_n_1634, mul_34_17_n_1635,
     mul_34_17_n_1636, mul_34_17_n_1637, mul_34_17_n_1638, mul_34_17_n_1639,
     mul_34_17_n_1640, mul_34_17_n_1641, mul_34_17_n_1642, mul_34_17_n_1643,
     mul_34_17_n_1644, mul_34_17_n_1645, mul_34_17_n_1646, mul_34_17_n_1647,
     mul_34_17_n_1648, mul_34_17_n_1649, mul_34_17_n_1650, mul_34_17_n_1651,
     mul_34_17_n_1652, mul_34_17_n_1653, mul_34_17_n_1654, mul_34_17_n_1655,
     mul_34_17_n_1656, mul_34_17_n_1657, mul_34_17_n_1658, mul_34_17_n_1659,
     mul_34_17_n_1660, mul_34_17_n_1661, mul_34_17_n_1662, mul_34_17_n_1663,
     mul_34_17_n_1664, mul_34_17_n_1665, mul_34_17_n_1666, mul_34_17_n_1667,
     mul_34_17_n_1668, mul_34_17_n_1669, mul_34_17_n_1670, mul_34_17_n_1671,
     mul_34_17_n_1672, mul_34_17_n_1673, mul_34_17_n_1674, mul_34_17_n_1675,
     mul_34_17_n_1676, mul_34_17_n_1677, mul_34_17_n_1678, mul_34_17_n_1679,
     mul_34_17_n_1680, mul_34_17_n_1681, mul_34_17_n_1682, mul_34_17_n_1683,
     mul_34_17_n_1684, mul_34_17_n_1685, mul_34_17_n_1686, mul_34_17_n_1687,
     mul_34_17_n_1688, mul_34_17_n_1689, mul_34_17_n_1690, mul_34_17_n_1691,
     mul_34_17_n_1692, mul_34_17_n_1693, mul_34_17_n_1694, mul_34_17_n_1695,
     mul_34_17_n_1696, mul_34_17_n_1697, mul_34_17_n_1698, mul_34_17_n_1699,
     mul_34_17_n_1700, mul_34_17_n_1701, mul_34_17_n_1702, mul_34_17_n_1703,
     mul_34_17_n_1704, mul_34_17_n_1705, mul_34_17_n_1706, mul_34_17_n_1707,
     mul_34_17_n_1708, mul_34_17_n_1709, mul_34_17_n_1710, mul_34_17_n_1711,
     mul_34_17_n_1712, mul_34_17_n_1713, mul_34_17_n_1714, mul_34_17_n_1715,
     mul_34_17_n_1716, mul_34_17_n_1717, mul_34_17_n_1718, mul_34_17_n_1719,
     mul_34_17_n_1720, mul_34_17_n_1721, mul_34_17_n_1722, mul_34_17_n_1723,
     mul_34_17_n_1724, mul_34_17_n_1725, mul_34_17_n_1726, mul_34_17_n_1727,
     mul_34_17_n_1728, mul_34_17_n_1729, mul_34_17_n_1730, mul_34_17_n_1731,
     mul_34_17_n_1732, mul_34_17_n_1733, mul_34_17_n_1734, mul_34_17_n_1735,
     mul_34_17_n_1736, mul_34_17_n_1737, mul_34_17_n_1738, mul_34_17_n_1739,
     mul_34_17_n_1740, mul_34_17_n_1741, mul_34_17_n_1742, mul_34_17_n_1743,
     mul_34_17_n_1744, mul_34_17_n_1745, mul_34_17_n_1746, mul_34_17_n_1747,
     mul_34_17_n_1748, mul_34_17_n_1749, mul_34_17_n_1750, mul_34_17_n_1751,
     mul_34_17_n_1752, mul_34_17_n_1753, mul_34_17_n_1754, mul_34_17_n_1755,
     mul_34_17_n_1756, mul_34_17_n_1757, mul_34_17_n_1758, mul_34_17_n_1759,
     mul_34_17_n_1760, mul_34_17_n_1761, mul_34_17_n_1762, mul_34_17_n_1763,
     mul_34_17_n_1764, mul_34_17_n_1765, mul_34_17_n_1766, mul_34_17_n_1767,
     mul_34_17_n_1768, mul_34_17_n_1769, mul_34_17_n_1770, mul_34_17_n_1771,
     mul_34_17_n_1772, mul_34_17_n_1773, mul_34_17_n_1774, mul_34_17_n_1775,
     mul_34_17_n_1776, mul_34_17_n_1777, mul_34_17_n_1778, mul_34_17_n_1779,
     mul_34_17_n_1780, mul_34_17_n_1781, mul_34_17_n_1782, mul_34_17_n_1783,
     mul_34_17_n_1784, mul_34_17_n_1785, mul_34_17_n_1786, mul_34_17_n_1787,
     mul_34_17_n_1788, mul_34_17_n_1789, mul_34_17_n_1790, mul_34_17_n_1791,
     mul_34_17_n_1792, mul_34_17_n_1793, mul_34_17_n_1794, mul_34_17_n_1795,
     mul_34_17_n_1796, mul_34_17_n_1797, mul_34_17_n_1798, mul_34_17_n_1799,
     mul_34_17_n_1800, mul_34_17_n_1801, mul_34_17_n_1802, mul_34_17_n_1803,
     mul_34_17_n_1804, mul_34_17_n_1805, mul_34_17_n_1806, mul_34_17_n_1807,
     mul_34_17_n_1808, mul_34_17_n_1809, mul_34_17_n_1810, mul_34_17_n_1811,
     mul_34_17_n_1812, mul_34_17_n_1813, mul_34_17_n_1814, mul_34_17_n_1815,
     mul_34_17_n_1816, mul_34_17_n_1817, mul_34_17_n_1818, mul_34_17_n_1819,
     mul_34_17_n_1820, mul_34_17_n_1821, mul_34_17_n_1822, mul_34_17_n_1823,
     mul_34_17_n_1824, mul_34_17_n_1825, mul_34_17_n_1826, mul_34_17_n_1827,
     mul_34_17_n_1828, mul_34_17_n_1829, mul_34_17_n_1830, mul_34_17_n_1831,
     mul_34_17_n_1832, mul_34_17_n_1833, mul_34_17_n_1834, mul_34_17_n_1835,
     mul_34_17_n_1836, mul_34_17_n_1837, mul_34_17_n_1838, mul_34_17_n_1839,
     mul_34_17_n_1840, mul_34_17_n_1841, mul_34_17_n_1842, mul_34_17_n_1843,
     mul_34_17_n_1844, mul_34_17_n_1845, mul_34_17_n_1846, mul_34_17_n_1847,
     mul_34_17_n_1848, mul_34_17_n_1849, mul_34_17_n_1850, mul_34_17_n_1851,
     mul_34_17_n_1852, mul_34_17_n_1853, mul_34_17_n_1854, mul_34_17_n_1855,
     mul_34_17_n_1856, mul_34_17_n_1857, mul_34_17_n_1858, mul_34_17_n_1859,
     mul_34_17_n_1860, mul_34_17_n_1861, mul_34_17_n_1862, mul_34_17_n_1863,
     mul_34_17_n_1864, mul_34_17_n_1865, mul_34_17_n_1866, mul_34_17_n_1867,
     mul_34_17_n_1868, mul_34_17_n_1869, mul_34_17_n_1870, mul_34_17_n_1871,
     mul_34_17_n_1872, mul_34_17_n_1873, mul_34_17_n_1874, mul_34_17_n_1875,
     mul_34_17_n_1876, mul_34_17_n_1877, mul_34_17_n_1878, mul_34_17_n_1879,
     mul_34_17_n_1880, mul_34_17_n_1881, mul_34_17_n_1882, mul_34_17_n_1883,
     mul_34_17_n_1884, mul_34_17_n_1885, mul_34_17_n_1886, mul_34_17_n_1887,
     mul_34_17_n_1888, mul_34_17_n_1889, mul_34_17_n_1890, mul_34_17_n_1891,
     mul_34_17_n_1892, mul_34_17_n_1893, mul_34_17_n_1894, mul_34_17_n_1895,
     mul_34_17_n_1896, mul_34_17_n_1897, mul_34_17_n_1898, mul_34_17_n_1899,
     mul_34_17_n_1900, mul_34_17_n_1901, mul_34_17_n_1902, mul_34_17_n_1903,
     mul_34_17_n_1904, mul_34_17_n_1905, mul_34_17_n_1906, mul_34_17_n_1907,
     mul_34_17_n_1908, mul_34_17_n_1909, mul_34_17_n_1910, mul_34_17_n_1911,
     mul_34_17_n_1912, mul_34_17_n_1913, mul_34_17_n_1914, mul_34_17_n_1915,
     mul_34_17_n_1916, mul_34_17_n_1917, mul_34_17_n_1918, mul_34_17_n_1919,
     mul_34_17_n_1920, mul_34_17_n_1921, mul_34_17_n_1922, mul_34_17_n_1923,
     mul_34_17_n_1924, mul_34_17_n_1925, mul_34_17_n_1926, mul_34_17_n_1927,
     mul_34_17_n_1928, mul_34_17_n_1929, mul_34_17_n_1930, mul_34_17_n_1931,
     mul_34_17_n_1932, mul_34_17_n_1933, mul_34_17_n_1934, mul_34_17_n_1935,
     mul_34_17_n_1936, mul_34_17_n_1937, mul_34_17_n_1938, mul_34_17_n_1939,
     mul_34_17_n_1940, mul_34_17_n_1941, mul_34_17_n_1942, mul_34_17_n_1943,
     mul_34_17_n_1944, mul_34_17_n_1945, mul_34_17_n_1946, mul_34_17_n_1947,
     mul_34_17_n_1948, mul_34_17_n_1949, mul_34_17_n_1950, mul_34_17_n_1951,
     mul_34_17_n_1952, mul_34_17_n_1953, mul_34_17_n_1954, mul_34_17_n_1955,
     mul_34_17_n_1956, mul_34_17_n_1957, mul_34_17_n_1958, mul_34_17_n_1959,
     mul_34_17_n_1960, mul_34_17_n_1961, mul_34_17_n_1962, mul_34_17_n_1963,
     mul_34_17_n_1964, mul_34_17_n_1965, mul_34_17_n_1966, mul_34_17_n_1967,
     mul_34_17_n_1968, mul_34_17_n_1969, mul_34_17_n_1970, mul_34_17_n_1971,
     mul_34_17_n_1972, mul_34_17_n_1973, mul_34_17_n_1974, mul_34_17_n_1975,
     mul_34_17_n_1976, mul_34_17_n_1977, mul_34_17_n_1978, mul_34_17_n_1979,
     mul_34_17_n_1980, mul_34_17_n_1981, mul_34_17_n_1982, mul_34_17_n_1983,
     mul_34_17_n_1984, mul_34_17_n_1985, mul_34_17_n_1986, mul_34_17_n_1987,
     mul_34_17_n_1988, mul_34_17_n_1989, mul_34_17_n_1990, mul_34_17_n_1991,
     mul_34_17_n_1992, mul_34_17_n_1993, mul_34_17_n_1994, mul_34_17_n_1995,
     mul_34_17_n_1996, mul_34_17_n_1997, mul_34_17_n_1998, mul_34_17_n_1999,
     mul_34_17_n_2000, mul_34_17_n_2001, mul_34_17_n_2002, mul_34_17_n_2003,
     mul_34_17_n_2004, mul_34_17_n_2005, mul_34_17_n_2006, mul_34_17_n_2007,
     mul_34_17_n_2008, mul_34_17_n_2009, mul_34_17_n_2010, mul_34_17_n_2011,
     mul_34_17_n_2012, mul_34_17_n_2013, mul_34_17_n_2014, mul_34_17_n_2015,
     mul_34_17_n_2016, mul_34_17_n_2017, mul_34_17_n_2018, mul_34_17_n_2019,
     mul_34_17_n_2020, mul_34_17_n_2021, mul_34_17_n_2022, mul_34_17_n_2023,
     mul_34_17_n_2024, mul_34_17_n_2025, mul_34_17_n_2026, mul_34_17_n_2027,
     mul_34_17_n_2028, mul_34_17_n_2029, mul_34_17_n_2030, mul_34_17_n_2031,
     mul_34_17_n_2032, mul_34_17_n_2033, mul_34_17_n_2034, mul_34_17_n_2035,
     mul_34_17_n_2036, mul_34_17_n_2037, mul_34_17_n_2038, mul_34_17_n_2039,
     mul_34_17_n_2040, mul_34_17_n_2041, mul_34_17_n_2042, mul_34_17_n_2043,
     mul_34_17_n_2044, mul_34_17_n_2045, mul_34_17_n_2046, mul_34_17_n_2047,
     mul_34_17_n_2048, mul_34_17_n_2049, mul_34_17_n_2050, mul_34_17_n_2051,
     mul_34_17_n_2052, mul_34_17_n_2053, mul_34_17_n_2054, mul_34_17_n_2055,
     mul_34_17_n_2056, mul_34_17_n_2057, mul_34_17_n_2058, mul_34_17_n_2059,
     mul_34_17_n_2060, mul_34_17_n_2061, mul_34_17_n_2062, mul_34_17_n_2063,
     mul_34_17_n_2064, mul_34_17_n_2065, mul_34_17_n_2066, mul_34_17_n_2067,
     mul_34_17_n_2068, mul_34_17_n_2069, mul_34_17_n_2070, mul_34_17_n_2071,
     mul_34_17_n_2072, mul_34_17_n_2073, mul_34_17_n_2074, mul_34_17_n_2075,
     mul_34_17_n_2076, mul_34_17_n_2077, mul_34_17_n_2078, mul_34_17_n_2079,
     mul_34_17_n_2080, mul_34_17_n_2081, mul_34_17_n_2082, mul_34_17_n_2083,
     mul_34_17_n_2084, mul_34_17_n_2085, mul_34_17_n_2086, mul_34_17_n_2087,
     mul_34_17_n_2088, mul_34_17_n_2089, mul_34_17_n_2090, mul_34_17_n_2091,
     mul_34_17_n_2092, mul_34_17_n_2093, mul_34_17_n_2094, mul_34_17_n_2095,
     mul_34_17_n_2096, mul_34_17_n_2097, mul_34_17_n_2098, mul_34_17_n_2099,
     mul_34_17_n_2100, mul_34_17_n_2101, mul_34_17_n_2102, mul_34_17_n_2103,
     mul_34_17_n_2104, mul_34_17_n_2105, mul_34_17_n_2106, mul_34_17_n_2107,
     mul_34_17_n_2108, mul_34_17_n_2109, mul_34_17_n_2110, mul_34_17_n_2111,
     mul_34_17_n_2112, mul_34_17_n_2113, mul_34_17_n_2114, mul_34_17_n_2115,
     mul_34_17_n_2116, mul_34_17_n_2117, mul_34_17_n_2118, mul_34_17_n_2119,
     mul_34_17_n_2120, mul_34_17_n_2121, mul_34_17_n_2122, mul_34_17_n_2123,
     mul_34_17_n_2124, mul_34_17_n_2125, mul_34_17_n_2126, mul_34_17_n_2127,
     mul_34_17_n_2128, mul_34_17_n_2129, mul_34_17_n_2130, mul_34_17_n_2131,
     mul_34_17_n_2132, mul_34_17_n_2133, mul_34_17_n_2134, mul_34_17_n_2135,
     mul_34_17_n_2136, mul_34_17_n_2137, mul_34_17_n_2138, mul_34_17_n_2139,
     mul_34_17_n_2140, mul_34_17_n_2141, mul_34_17_n_2142, mul_34_17_n_2143,
     mul_34_17_n_2144, mul_34_17_n_2145, mul_34_17_n_2146, mul_34_17_n_2147,
     mul_34_17_n_2148, mul_34_17_n_2149, mul_34_17_n_2150, mul_34_17_n_2151,
     mul_34_17_n_2152, mul_34_17_n_2153, mul_34_17_n_2154, mul_34_17_n_2155,
     mul_34_17_n_2156, mul_34_17_n_2157, mul_34_17_n_2158, mul_34_17_n_2159,
     mul_34_17_n_2160, mul_34_17_n_2161, mul_34_17_n_2162, mul_34_17_n_2163,
     mul_34_17_n_2164, mul_34_17_n_2165, mul_34_17_n_2166, mul_34_17_n_2167,
     mul_34_17_n_2168, mul_34_17_n_2169, mul_34_17_n_2170, mul_34_17_n_2171,
     mul_34_17_n_2172, mul_34_17_n_2173, mul_34_17_n_2174, mul_34_17_n_2175,
     mul_34_17_n_2176, mul_34_17_n_2177, mul_34_17_n_2178, mul_34_17_n_2179,
     mul_34_17_n_2180, mul_34_17_n_2181, mul_34_17_n_2182, mul_34_17_n_2183,
     mul_34_17_n_2184, mul_34_17_n_2185, mul_34_17_n_2186, mul_34_17_n_2187,
     mul_34_17_n_2188, mul_34_17_n_2189, mul_34_17_n_2190, mul_34_17_n_2191,
     mul_34_17_n_2192, mul_34_17_n_2193, mul_34_17_n_2194, mul_34_17_n_2195,
     mul_34_17_n_2196, mul_34_17_n_2197, mul_34_17_n_2198, mul_34_17_n_2199,
     mul_34_17_n_2200, mul_34_17_n_2201, mul_34_17_n_2202, mul_34_17_n_2203,
     mul_34_17_n_2204, mul_34_17_n_2205, mul_34_17_n_2206, mul_34_17_n_2207,
     mul_34_17_n_2208, mul_34_17_n_2209, mul_34_17_n_2210, mul_34_17_n_2211,
     mul_34_17_n_2212, mul_34_17_n_2213, mul_34_17_n_2214, mul_34_17_n_2215,
     mul_34_17_n_2216, mul_34_17_n_2217, mul_34_17_n_2218, mul_34_17_n_2219,
     mul_34_17_n_2220, mul_34_17_n_2221, mul_34_17_n_2222, mul_34_17_n_2223,
     mul_34_17_n_2224, mul_34_17_n_2225, mul_34_17_n_2226, mul_34_17_n_2227,
     mul_34_17_n_2228, mul_34_17_n_2229, mul_34_17_n_2230, mul_34_17_n_2231,
     mul_34_17_n_2232, mul_34_17_n_2233, mul_34_17_n_2234, mul_34_17_n_2235,
     mul_34_17_n_2236, mul_34_17_n_2237, mul_34_17_n_2238, mul_34_17_n_2239,
     mul_34_17_n_2240, mul_34_17_n_2241, mul_34_17_n_2242, mul_34_17_n_2243,
     mul_34_17_n_2244, mul_34_17_n_2245, mul_34_17_n_2246, mul_34_17_n_2247,
     mul_34_17_n_2248, mul_34_17_n_2249, mul_34_17_n_2250, mul_34_17_n_2251,
     mul_34_17_n_2252, mul_34_17_n_2253, mul_34_17_n_2254, mul_34_17_n_2255,
     mul_34_17_n_2256, mul_34_17_n_2257, mul_34_17_n_2258, mul_34_17_n_2259,
     mul_34_17_n_2260, mul_34_17_n_2261, mul_34_17_n_2262, mul_34_17_n_2263,
     mul_34_17_n_2264, mul_34_17_n_2265, mul_34_17_n_2266, mul_34_17_n_2267,
     mul_34_17_n_2268, mul_34_17_n_2269, mul_34_17_n_2270, mul_34_17_n_2271,
     mul_34_17_n_2272, mul_34_17_n_2273, mul_34_17_n_2274, mul_34_17_n_2275,
     mul_34_17_n_2276, mul_34_17_n_2277, mul_34_17_n_2278, mul_34_17_n_2279,
     mul_34_17_n_2280, mul_34_17_n_2281, mul_34_17_n_2282, mul_34_17_n_2283,
     mul_34_17_n_2284, mul_34_17_n_2285, mul_34_17_n_2286, mul_34_17_n_2287,
     mul_34_17_n_2288, mul_34_17_n_2289, mul_34_17_n_2290, mul_34_17_n_2291,
     mul_34_17_n_2292, mul_34_17_n_2293, mul_34_17_n_2294, mul_34_17_n_2295,
     mul_34_17_n_2296, mul_34_17_n_2297, mul_34_17_n_2298, mul_34_17_n_2299,
     mul_34_17_n_2300, mul_34_17_n_2301, mul_34_17_n_2302, mul_34_17_n_2303,
     mul_34_17_n_2304, mul_34_17_n_2305, mul_34_17_n_2306, mul_34_17_n_2307,
     mul_34_17_n_2308, mul_34_17_n_2309, mul_34_17_n_2310, mul_34_17_n_2311,
     mul_34_17_n_2312, mul_34_17_n_2313, mul_34_17_n_2314, mul_34_17_n_2315,
     mul_34_17_n_2316, mul_34_17_n_2317, mul_34_17_n_2318, mul_34_17_n_2319,
     mul_34_17_n_2320, mul_34_17_n_2321, mul_34_17_n_2322, mul_34_17_n_2323,
     mul_34_17_n_2324, mul_34_17_n_2325, mul_34_17_n_2326, mul_34_17_n_2327,
     mul_34_17_n_2328, mul_34_17_n_2329, mul_34_17_n_2330, mul_34_17_n_2331,
     mul_34_17_n_2332, mul_34_17_n_2333, mul_34_17_n_2334, mul_34_17_n_2335,
     mul_34_17_n_2336, mul_34_17_n_2337, mul_34_17_n_2338, mul_34_17_n_2339,
     mul_34_17_n_2340, mul_34_17_n_2341, mul_34_17_n_2342, mul_34_17_n_2343,
     mul_34_17_n_2344, mul_34_17_n_2345, mul_34_17_n_2346, mul_34_17_n_2347,
     mul_34_17_n_2348, mul_34_17_n_2349, mul_34_17_n_2350, mul_34_17_n_2351,
     mul_34_17_n_2352, mul_34_17_n_2353, mul_34_17_n_2354, mul_34_17_n_2355,
     mul_34_17_n_2356, mul_34_17_n_2357, mul_34_17_n_2358, mul_34_17_n_2359,
     mul_34_17_n_2360, mul_34_17_n_2361, mul_34_17_n_2362, mul_34_17_n_2363,
     mul_34_17_n_2364, mul_34_17_n_2365, mul_34_17_n_2366, mul_34_17_n_2367,
     mul_34_17_n_2368, mul_34_17_n_2369, mul_34_17_n_2370, mul_34_17_n_2371,
     mul_34_17_n_2372, mul_34_17_n_2373, mul_34_17_n_2374, mul_34_17_n_2375,
     mul_34_17_n_2376, mul_34_17_n_2377, mul_34_17_n_2378, mul_34_17_n_2379,
     mul_34_17_n_2380, mul_34_17_n_2381, mul_34_17_n_2382, mul_34_17_n_2383,
     mul_34_17_n_2384, mul_34_17_n_2385, mul_34_17_n_2386, mul_34_17_n_2387,
     mul_34_17_n_2388, mul_34_17_n_2389, mul_34_17_n_2390, mul_34_17_n_2391,
     mul_34_17_n_2392, mul_34_17_n_2393, mul_34_17_n_2394, mul_34_17_n_2395,
     mul_34_17_n_2396, mul_34_17_n_2397, mul_34_17_n_2398, mul_34_17_n_2399,
     mul_34_17_n_2400, mul_34_17_n_2401, mul_34_17_n_2402, mul_34_17_n_2403,
     mul_34_17_n_2404, mul_34_17_n_2405, mul_34_17_n_2406, mul_34_17_n_2407,
     mul_34_17_n_2408, mul_34_17_n_2409, mul_34_17_n_2410, mul_34_17_n_2411,
     mul_34_17_n_2412, mul_34_17_n_2413, mul_34_17_n_2414, mul_34_17_n_2415,
     mul_34_17_n_2416, mul_34_17_n_2417, mul_34_17_n_2418, mul_34_17_n_2419,
     mul_34_17_n_2420, mul_34_17_n_2421, mul_34_17_n_2422, mul_34_17_n_2423,
     mul_34_17_n_2424, mul_34_17_n_2425, mul_34_17_n_2426, mul_34_17_n_2427,
     mul_34_17_n_2428, mul_34_17_n_2429, mul_34_17_n_2430, mul_34_17_n_2431,
     mul_34_17_n_2432, mul_34_17_n_2433, mul_34_17_n_2434, mul_34_17_n_2435,
     mul_34_17_n_2436, mul_34_17_n_2437, mul_34_17_n_2438, mul_34_17_n_2439,
     mul_34_17_n_2440, mul_34_17_n_2441, mul_34_17_n_2442, mul_34_17_n_2443,
     mul_34_17_n_2444, mul_34_17_n_2445, mul_34_17_n_2446, mul_34_17_n_2447,
     mul_34_17_n_2448, mul_34_17_n_2449, mul_34_17_n_2450, mul_34_17_n_2451,
     mul_34_17_n_2452, mul_34_17_n_2453, mul_34_17_n_2454, mul_34_17_n_2455,
     mul_34_17_n_2456, mul_34_17_n_2457, mul_34_17_n_2458, mul_34_17_n_2459,
     mul_34_17_n_2460, mul_34_17_n_2461, mul_34_17_n_2462, mul_34_17_n_2463,
     mul_34_17_n_2464, mul_34_17_n_2465, mul_34_17_n_2466, mul_34_17_n_2467,
     mul_34_17_n_2468, mul_34_17_n_2469, mul_34_17_n_2470, mul_34_17_n_2471,
     mul_34_17_n_2472, mul_34_17_n_2473, mul_34_17_n_2474, mul_34_17_n_2475,
     mul_34_17_n_2476, mul_34_17_n_2477, mul_34_17_n_2478, mul_34_17_n_2479,
     mul_34_17_n_2480, mul_34_17_n_2481, mul_34_17_n_2482, mul_34_17_n_2483,
     mul_34_17_n_2484, mul_34_17_n_2485, mul_34_17_n_2486, mul_34_17_n_2487,
     mul_34_17_n_2488, mul_34_17_n_2489, mul_34_17_n_2490, mul_34_17_n_2491,
     mul_34_17_n_2492, mul_34_17_n_2493, mul_34_17_n_2494, mul_34_17_n_2495,
     mul_34_17_n_2496, mul_34_17_n_2497, mul_34_17_n_2498, mul_34_17_n_2499,
     mul_34_17_n_2500, mul_34_17_n_2501, mul_34_17_n_2502, mul_34_17_n_2503,
     mul_34_17_n_2504, mul_34_17_n_2505, mul_34_17_n_2506, mul_34_17_n_2507,
     mul_34_17_n_2508, mul_34_17_n_2509, mul_34_17_n_2510, mul_34_17_n_2511,
     mul_34_17_n_2512, mul_34_17_n_2513, mul_34_17_n_2514, mul_34_17_n_2515,
     mul_34_17_n_2516, mul_34_17_n_2517, mul_34_17_n_2518, mul_34_17_n_2519,
     mul_34_17_n_2520, mul_34_17_n_2521, mul_34_17_n_2522, mul_34_17_n_2523,
     mul_34_17_n_2524, mul_34_17_n_2525, mul_34_17_n_2526, mul_34_17_n_2527,
     mul_34_17_n_2528, mul_34_17_n_2529, mul_34_17_n_2530, mul_34_17_n_2531,
     mul_34_17_n_2532, mul_34_17_n_2533, mul_34_17_n_2534, mul_34_17_n_2535,
     mul_34_17_n_2536, mul_34_17_n_2537, mul_34_17_n_2538, mul_34_17_n_2539,
     mul_34_17_n_2540, mul_34_17_n_2541, mul_34_17_n_2542, mul_34_17_n_2543,
     mul_34_17_n_2544, mul_34_17_n_2545, mul_34_17_n_2546, mul_34_17_n_2547,
     mul_34_17_n_2548, mul_34_17_n_2549, mul_34_17_n_2550, mul_34_17_n_2551,
     mul_34_17_n_2552, mul_34_17_n_2553, mul_34_17_n_2554, mul_34_17_n_2555,
     mul_34_17_n_2556, mul_34_17_n_2557, mul_34_17_n_2558, mul_34_17_n_2559,
     mul_34_17_n_2560, mul_34_17_n_2561, mul_34_17_n_2562, mul_34_17_n_2563,
     mul_34_17_n_2564, mul_34_17_n_2565, mul_34_17_n_2566, mul_34_17_n_2567,
     mul_34_17_n_2568, mul_34_17_n_2569, mul_34_17_n_2570, mul_34_17_n_2571,
     mul_34_17_n_2572, mul_34_17_n_2573, mul_34_17_n_2574, mul_34_17_n_2575,
     mul_34_17_n_2576, mul_34_17_n_2577, mul_34_17_n_2578, mul_34_17_n_2579,
     mul_34_17_n_2580, mul_34_17_n_2581, mul_34_17_n_2582, mul_34_17_n_2583,
     mul_34_17_n_2584, mul_34_17_n_2585, mul_34_17_n_2586, mul_34_17_n_2587,
     mul_34_17_n_2588, mul_34_17_n_2589, mul_34_17_n_2590, mul_34_17_n_2591,
     mul_34_17_n_2592, mul_34_17_n_2593, mul_34_17_n_2594, mul_34_17_n_2595,
     mul_34_17_n_2596, mul_34_17_n_2597, mul_34_17_n_2598, mul_34_17_n_2599,
     mul_34_17_n_2600, mul_34_17_n_2601, mul_34_17_n_2602, mul_34_17_n_2603,
     mul_34_17_n_2604, mul_34_17_n_2605, mul_34_17_n_2606, mul_34_17_n_2607,
     mul_34_17_n_2608, mul_34_17_n_2609, mul_34_17_n_2610, mul_34_17_n_2611,
     mul_34_17_n_2612, mul_34_17_n_2613, mul_34_17_n_2614, mul_34_17_n_2615,
     mul_34_17_n_2616, mul_34_17_n_2617, mul_34_17_n_2618, mul_34_17_n_2619,
     mul_34_17_n_2620, mul_34_17_n_2621, mul_34_17_n_2622, mul_34_17_n_2623,
     mul_34_17_n_2624, mul_34_17_n_2625, mul_34_17_n_2626, mul_34_17_n_2627,
     mul_34_17_n_2628, mul_34_17_n_2629, mul_34_17_n_2630, mul_34_17_n_2631,
     mul_34_17_n_2632, mul_34_17_n_2633, mul_34_17_n_2634, mul_34_17_n_2635,
     mul_34_17_n_2636, mul_34_17_n_2637, mul_34_17_n_2638, mul_34_17_n_2639,
     mul_34_17_n_2640, mul_34_17_n_2641, mul_34_17_n_2642, mul_34_17_n_2643,
     mul_34_17_n_2644, mul_34_17_n_2645, mul_34_17_n_2646, mul_34_17_n_2647,
     mul_34_17_n_2648, mul_34_17_n_2649, mul_34_17_n_2650, mul_34_17_n_2651,
     mul_34_17_n_2652, mul_34_17_n_2653, mul_34_17_n_2654, mul_34_17_n_2655,
     mul_34_17_n_2656, mul_34_17_n_2657, mul_34_17_n_2658, mul_34_17_n_2659,
     mul_34_17_n_2660, mul_34_17_n_2661, mul_34_17_n_2662, mul_34_17_n_2663,
     mul_34_17_n_2664, mul_34_17_n_2665, mul_34_17_n_2666, mul_34_17_n_2667,
     mul_34_17_n_2668, mul_34_17_n_2669, mul_34_17_n_2670, mul_34_17_n_2671,
     mul_34_17_n_2672, mul_34_17_n_2673, mul_34_17_n_2674, mul_34_17_n_2675,
     mul_34_17_n_2676, mul_34_17_n_2677, mul_34_17_n_2678, mul_34_17_n_2679,
     mul_34_17_n_2680, mul_34_17_n_2681, mul_34_17_n_2682, mul_34_17_n_2683,
     mul_34_17_n_2684, mul_34_17_n_2685, mul_34_17_n_2686, mul_34_17_n_2687,
     mul_34_17_n_2688, mul_34_17_n_2689, mul_34_17_n_2690, mul_34_17_n_2691,
     mul_34_17_n_2692, mul_34_17_n_2693, mul_34_17_n_2694, mul_34_17_n_2695,
     mul_34_17_n_2696, mul_34_17_n_2697, mul_34_17_n_2698, mul_34_17_n_2699,
     mul_34_17_n_2700, mul_34_17_n_2701, mul_34_17_n_2702, mul_34_17_n_2703,
     mul_34_17_n_2704, mul_34_17_n_2705, mul_34_17_n_2706, mul_34_17_n_2707,
     mul_34_17_n_2708, mul_34_17_n_2709, mul_34_17_n_2710, mul_34_17_n_2711,
     mul_34_17_n_2712, mul_34_17_n_2713, mul_34_17_n_2714, mul_34_17_n_2715,
     mul_34_17_n_2716, mul_34_17_n_2717, mul_34_17_n_2718, mul_34_17_n_2719,
     mul_34_17_n_2720, mul_34_17_n_2721, mul_34_17_n_2722, mul_34_17_n_2723,
     mul_34_17_n_2724, mul_34_17_n_2725, mul_34_17_n_2726, mul_34_17_n_2727,
     mul_34_17_n_2728, mul_34_17_n_2729, mul_34_17_n_2730, mul_34_17_n_2731,
     mul_34_17_n_2732, mul_34_17_n_2733, mul_34_17_n_2734, mul_34_17_n_2735,
     mul_34_17_n_2736, mul_34_17_n_2737, mul_34_17_n_2738, mul_34_17_n_2739,
     mul_34_17_n_2740, mul_34_17_n_2741, mul_34_17_n_2742, mul_34_17_n_2743,
     mul_34_17_n_2744, mul_34_17_n_2745, mul_34_17_n_2746, mul_34_17_n_2747,
     mul_34_17_n_2748, mul_34_17_n_2749, mul_34_17_n_2750, mul_34_17_n_2751,
     mul_34_17_n_2752, mul_34_17_n_2753, mul_34_17_n_2754, mul_34_17_n_2755,
     mul_34_17_n_2756, mul_34_17_n_2757, mul_34_17_n_2758, mul_34_17_n_2759,
     mul_34_17_n_2760, mul_34_17_n_2761, mul_34_17_n_2762, mul_34_17_n_2763,
     mul_34_17_n_2764, mul_34_17_n_2765, mul_34_17_n_2766, mul_34_17_n_2767,
     mul_34_17_n_2768, mul_34_17_n_2769, mul_34_17_n_2770, mul_34_17_n_2771,
     mul_34_17_n_2772, mul_34_17_n_2773, mul_34_17_n_2774, mul_34_17_n_2775,
     mul_34_17_n_2776, mul_34_17_n_2777, mul_34_17_n_2809, mul_34_17_n_2810,
     mul_34_17_n_2811, mul_34_17_n_2812, mul_34_17_n_2813, mul_34_17_n_2814,
     mul_34_17_n_2815, mul_34_17_n_2816, mul_34_17_n_2817, mul_34_17_n_2818,
     mul_34_17_n_2819, mul_34_17_n_2820, mul_34_17_n_2821, mul_34_17_n_2822,
     mul_34_17_n_2823, mul_34_17_n_2824, mul_34_17_n_2825, mul_34_17_n_2826,
     mul_34_17_n_2827, mul_34_17_n_2828, mul_34_17_n_2829, mul_34_17_n_2830,
     mul_34_17_n_2831, mul_34_17_n_2832, mul_34_17_n_2833, mul_34_17_n_2834,
     mul_34_17_n_2835, mul_34_17_n_2836, mul_34_17_n_2837, mul_34_17_n_2838,
     mul_34_17_n_2839, mul_34_17_n_2840, mul_34_17_n_2841, mul_34_17_n_2842,
     mul_34_17_n_2843, mul_34_17_n_2844, mul_34_17_n_2845, mul_34_17_n_2846,
     mul_34_17_n_2847, mul_34_17_n_2848, mul_34_17_n_2849, mul_34_17_n_2850,
     mul_34_17_n_2851, mul_34_17_n_2852, mul_34_17_n_2853, mul_34_17_n_2854,
     mul_34_17_n_2855, mul_34_17_n_2856, mul_34_17_n_2857, mul_34_17_n_2858,
     mul_34_17_n_2859, mul_34_17_n_2860, mul_34_17_n_2861, mul_34_17_n_2862,
     mul_34_17_n_2863, mul_34_17_n_2864, mul_34_17_n_2865, mul_34_17_n_2866,
     mul_34_17_n_2867, mul_34_17_n_2868, mul_34_17_n_2869, mul_34_17_n_2870,
     mul_34_17_n_2871, mul_34_17_n_2872, mul_34_17_n_2873, mul_34_17_n_2874,
     mul_34_17_n_2875, mul_34_17_n_2876, mul_34_17_n_2877, mul_34_17_n_2878,
     mul_34_17_n_2880, mul_34_17_n_2882, mul_34_17_n_2884, mul_34_17_n_2886,
     mul_34_17_n_2888, mul_34_17_n_2890, mul_34_17_n_2894, mul_34_17_n_2896,
     mul_34_17_n_2898, mul_34_17_n_2900, mul_34_17_n_2902, mul_34_17_n_2904,
     mul_34_17_n_2906, mul_34_17_n_2908, mul_34_17_n_2910, mul_34_17_n_2912,
     mul_34_17_n_2914, mul_34_17_n_2916, mul_34_17_n_2918, mul_34_17_n_2920,
     mul_34_17_n_2922, mul_34_17_n_2924, mul_34_17_n_2926, mul_34_17_n_2928,
     mul_34_17_n_2931, mul_34_17_n_2933, mul_34_17_n_2936, mul_34_17_n_2938,
     mul_34_17_n_2939, mul_34_17_n_2940, mul_34_17_n_2941, mul_34_17_n_2942,
     mul_34_17_n_2943, mul_34_17_n_2944, mul_34_17_n_2945, mul_34_17_n_2946,
     mul_34_17_n_2947, mul_34_17_n_2948, mul_34_17_n_2949, mul_34_17_n_2950,
     mul_34_17_n_2951, mul_34_17_n_2952, mul_34_17_n_2953, mul_34_17_n_2954,
     mul_34_17_n_2955, mul_34_17_n_2956, mul_34_17_n_2957, mul_34_17_n_2958,
     mul_34_17_n_2959, mul_34_17_n_2960, mul_34_17_n_2961, mul_34_17_n_2962,
     mul_34_17_n_2963, mul_34_17_n_2964, mul_34_17_n_2965, mul_34_17_n_2966,
     mul_34_17_n_2967, mul_34_17_n_2968, mul_34_17_n_2969, mul_34_17_n_2970,
     mul_34_17_n_2972, mul_34_17_n_2973, mul_34_17_n_2974, mul_34_17_n_2975,
     mul_34_17_n_2976, mul_34_17_n_2977, mul_34_17_n_2978, mul_34_17_n_2979,
     mul_34_17_n_2980, mul_34_17_n_2981, mul_34_17_n_2982, mul_34_17_n_2983,
     mul_34_17_n_2984, mul_34_17_n_2985, mul_34_17_n_2986, mul_34_17_n_2987,
     mul_34_17_n_2988, mul_34_17_n_2989, mul_34_17_n_2990, mul_34_17_n_2992,
     mul_34_17_n_2993, mul_34_17_n_2994, mul_34_17_n_2995, mul_34_17_n_2996,
     mul_34_17_n_2997, mul_34_17_n_2998, mul_34_17_n_2999, mul_34_17_n_3000,
     mul_34_17_n_3001, mul_34_17_n_3002, mul_34_17_n_3003, mul_34_17_n_3004,
     mul_34_17_n_3005, mul_34_17_n_3006, mul_34_17_n_3007, mul_34_17_n_3008,
     mul_34_17_n_3009, mul_34_17_n_3010, mul_34_17_n_3011, mul_34_17_n_3012,
     mul_34_17_n_3013, mul_34_17_n_3014, mul_34_17_n_3015, mul_34_17_n_3016,
     mul_34_17_n_3017, mul_34_17_n_3018, mul_34_17_n_3019, mul_34_17_n_3020,
     mul_34_17_n_3021, mul_34_17_n_3022, mul_34_17_n_3023, mul_34_17_n_3024,
     mul_34_17_n_3025, mul_34_17_n_3026, mul_34_17_n_3027, mul_34_17_n_3028,
     mul_34_17_n_3029, mul_34_17_n_3030, mul_34_17_n_3031, mul_34_17_n_3032,
     mul_34_17_n_3033, mul_34_17_n_3034, mul_34_17_n_3035, mul_34_17_n_3036,
     mul_34_17_n_3037, mul_34_17_n_3038, mul_34_17_n_3039, mul_34_17_n_3040,
     mul_34_17_n_3041, mul_34_17_n_3042, mul_34_17_n_3043, mul_34_17_n_3044,
     mul_34_17_n_3045, mul_34_17_n_3046, mul_34_17_n_3047, mul_34_17_n_3048,
     mul_34_17_n_3049, mul_34_17_n_3050, mul_34_17_n_3051, mul_34_17_n_3052,
     mul_34_17_n_3053, mul_34_17_n_3054, mul_34_17_n_3055, mul_34_17_n_3056,
     mul_34_17_n_3057, mul_34_17_n_3058, mul_34_17_n_3059, mul_34_17_n_3060,
     mul_34_17_n_3061, mul_34_17_n_3062, mul_34_17_n_3063, mul_34_17_n_3064,
     mul_34_17_n_3065, mul_34_17_n_3066, mul_34_17_n_3067, mul_34_17_n_3068,
     mul_34_17_n_3069, mul_34_17_n_3070, mul_34_17_n_3071, mul_34_17_n_3072,
     mul_34_17_n_3073, mul_34_17_n_3074, mul_34_17_n_3075, mul_34_17_n_3076,
     mul_34_17_n_3077, mul_34_17_n_3078, mul_34_17_n_3079, mul_34_17_n_3080,
     mul_34_17_n_3081, mul_34_17_n_3082, mul_34_17_n_3083, mul_34_17_n_3084,
     mul_34_17_n_3085, mul_34_17_n_3086, mul_34_17_n_3087, mul_34_17_n_3088,
     mul_34_17_n_3089, mul_34_17_n_3090, mul_34_17_n_3091, mul_34_17_n_3092,
     mul_34_17_n_3093, mul_34_17_n_3094, mul_34_17_n_3095, mul_34_17_n_3096,
     mul_34_17_n_3097, mul_34_17_n_3098, mul_34_17_n_3099, mul_34_17_n_3100,
     mul_34_17_n_3101, mul_34_17_n_3102, mul_34_17_n_3103, mul_34_17_n_3104,
     mul_34_17_n_3105, mul_34_17_n_3106, mul_34_17_n_3107, mul_34_17_n_3108,
     mul_34_17_n_3109, mul_34_17_n_3110, mul_34_17_n_3111, mul_34_17_n_3112,
     mul_34_17_n_3113, mul_34_17_n_3114, mul_34_17_n_3115, mul_34_17_n_3116,
     mul_34_17_n_3117, mul_34_17_n_3118, mul_34_17_n_3119, mul_34_17_n_3120,
     mul_34_17_n_3121, mul_34_17_n_3122, mul_34_17_n_3123, mul_34_17_n_3124,
     mul_34_17_n_3125, mul_34_17_n_3126, mul_34_17_n_3127, mul_34_17_n_3128,
     mul_34_17_n_3129, mul_34_17_n_3130, mul_34_17_n_3131, mul_34_17_n_3132,
     mul_34_17_n_3133, mul_34_17_n_3134, mul_34_17_n_3135, mul_34_17_n_3136,
     mul_34_17_n_3137, mul_34_17_n_3138, mul_34_17_n_3139, mul_34_17_n_3140,
     mul_34_17_n_3141, mul_34_17_n_3142, mul_34_17_n_3143, mul_34_17_n_3144,
     mul_34_17_n_3145, mul_34_17_n_3146, mul_34_17_n_3147, mul_34_17_n_3148,
     mul_34_17_n_3149, mul_34_17_n_3150, mul_34_17_n_3151, mul_34_17_n_3152,
     mul_34_17_n_3153, mul_34_17_n_3154, mul_34_17_n_3155, mul_34_17_n_3156,
     mul_34_17_n_3157, mul_34_17_n_3158, mul_34_17_n_3159, mul_34_17_n_3160,
     mul_34_17_n_3161, mul_34_17_n_3162, mul_34_17_n_3163, mul_34_17_n_3164,
     mul_34_17_n_3165, mul_34_17_n_3166, mul_34_17_n_3167, mul_34_17_n_3168,
     mul_34_17_n_3169, mul_34_17_n_3170, mul_34_17_n_3171, mul_34_17_n_3172,
     mul_34_17_n_3173, mul_34_17_n_3174, mul_34_17_n_3175, mul_34_17_n_3176,
     mul_34_17_n_3177, mul_34_17_n_3178, mul_34_17_n_3179, mul_34_17_n_3180,
     mul_34_17_n_3181, mul_34_17_n_3182, mul_34_17_n_3183, mul_34_17_n_3184,
     mul_34_17_n_3185, mul_34_17_n_3186, mul_34_17_n_3187, mul_34_17_n_3188,
     mul_34_17_n_3189, mul_34_17_n_3190, mul_34_17_n_3191, mul_34_17_n_3192,
     mul_34_17_n_3193, mul_34_17_n_3194, mul_34_17_n_3195, mul_34_17_n_3196,
     mul_34_17_n_3197, mul_34_17_n_3198, mul_34_17_n_3199, mul_34_17_n_3200,
     mul_34_17_n_3201, mul_34_17_n_3202, mul_34_17_n_3203, mul_34_17_n_3204,
     mul_34_17_n_3205, mul_34_17_n_3206, mul_34_17_n_3207, mul_34_17_n_3208,
     mul_34_17_n_3209, mul_34_17_n_3210, mul_34_17_n_3211, mul_34_17_n_3212,
     mul_34_17_n_3213, mul_34_17_n_3214, mul_34_17_n_3215, mul_34_17_n_3216,
     mul_34_17_n_3217, mul_34_17_n_3218, mul_34_17_n_3219, mul_34_17_n_3220,
     mul_34_17_n_3221, mul_34_17_n_3222, mul_34_17_n_3223, mul_34_17_n_3224,
     mul_34_17_n_3225, mul_34_17_n_3226, mul_34_17_n_3227, mul_34_17_n_3228,
     mul_34_17_n_3229, mul_34_17_n_3230, mul_34_17_n_3231, mul_34_17_n_3232,
     mul_34_17_n_3234, mul_34_17_n_3235, mul_34_17_n_3236, mul_34_17_n_3237,
     mul_34_17_n_3238, mul_34_17_n_3239, mul_34_17_n_3240, mul_34_17_n_3241,
     mul_34_17_n_3242, mul_34_17_n_3243, mul_34_17_n_3244, mul_34_17_n_3245,
     mul_34_17_n_3246, mul_34_17_n_3247, mul_34_17_n_3248, mul_34_17_n_3249,
     mul_34_17_n_3250, mul_34_17_n_3251, mul_34_17_n_3252, mul_34_17_n_3253,
     mul_34_17_n_3254, mul_34_17_n_3255, mul_34_17_n_3256, mul_34_17_n_3257,
     mul_34_17_n_3258, mul_34_17_n_3259, mul_34_17_n_3260, mul_34_17_n_3261,
     mul_34_17_n_3262, mul_34_17_n_3263, mul_34_17_n_3264, mul_34_17_n_3265,
     mul_34_17_n_3266, mul_34_17_n_3267, mul_34_17_n_3268, mul_34_17_n_3269,
     mul_34_17_n_3270, mul_34_17_n_3271, mul_34_17_n_3272, mul_34_17_n_3273,
     mul_34_17_n_3274, mul_34_17_n_3275, mul_34_17_n_3276, mul_34_17_n_3277,
     mul_34_17_n_3278, mul_34_17_n_3279, mul_34_17_n_3280, mul_34_17_n_3281,
     mul_34_17_n_3282, mul_34_17_n_3283, mul_34_17_n_3284, mul_34_17_n_3285,
     mul_34_17_n_3286, mul_34_17_n_3287, mul_34_17_n_3288, mul_34_17_n_3289,
     mul_34_17_n_3290, mul_34_17_n_3291, mul_34_17_n_3292, mul_34_17_n_3293,
     mul_34_17_n_3294, mul_34_17_n_3295, mul_34_17_n_3296, mul_34_17_n_3297,
     mul_34_17_n_3298, mul_34_17_n_3299, mul_34_17_n_3300, mul_34_17_n_3301,
     mul_34_17_n_3302, mul_34_17_n_3303, mul_34_17_n_3304, mul_34_17_n_3305,
     mul_34_17_n_3306, mul_34_17_n_3307, mul_34_17_n_3308, mul_34_17_n_3309,
     mul_34_17_n_3310, mul_34_17_n_3311, mul_34_17_n_3312, mul_34_17_n_3313,
     mul_34_17_n_3314, mul_34_17_n_3315, mul_34_17_n_3316, mul_34_17_n_3317,
     mul_34_17_n_3318, mul_34_17_n_3319, mul_34_17_n_3320, mul_34_17_n_3321,
     mul_34_17_n_3322, mul_34_17_n_3323, mul_34_17_n_3324, mul_34_17_n_3325,
     mul_34_17_n_3326, mul_34_17_n_3327, mul_34_17_n_3328, mul_34_17_n_3329,
     mul_34_17_n_3330, mul_34_17_n_3331, mul_34_17_n_3332, mul_34_17_n_3333,
     mul_34_17_n_3334, mul_34_17_n_3335, mul_34_17_n_3336, mul_34_17_n_3337,
     mul_34_17_n_3338, mul_34_17_n_3339, mul_34_17_n_3340, mul_34_17_n_3341,
     mul_34_17_n_3342, mul_34_17_n_3343, mul_34_17_n_3344, mul_34_17_n_3345,
     mul_34_17_n_3346, mul_34_17_n_3347, mul_34_17_n_3348, mul_34_17_n_3349,
     mul_34_17_n_3350, mul_34_17_n_3351, mul_34_17_n_3352, mul_34_17_n_3353,
     mul_34_17_n_3354, mul_34_17_n_3355, mul_34_17_n_3356, mul_34_17_n_3357,
     mul_34_17_n_3358, mul_34_17_n_3359, mul_34_17_n_3360, mul_34_17_n_3361,
     mul_34_17_n_3362, mul_34_17_n_3363, mul_34_17_n_3364, mul_34_17_n_3365,
     mul_34_17_n_3366, mul_34_17_n_3367, mul_34_17_n_3368, mul_34_17_n_3369,
     mul_34_17_n_3370, mul_34_17_n_3371, mul_34_17_n_3372, mul_34_17_n_3373,
     mul_34_17_n_3374, mul_34_17_n_3375, mul_34_17_n_3376, mul_34_17_n_3377,
     mul_34_17_n_3378, mul_34_17_n_3379, mul_34_17_n_3380, mul_34_17_n_3381,
     mul_34_17_n_3382, mul_34_17_n_3383, mul_34_17_n_3384, mul_34_17_n_3385,
     mul_34_17_n_3386, mul_34_17_n_3387, mul_34_17_n_3388, mul_34_17_n_3389,
     mul_34_17_n_3390, mul_34_17_n_3391, mul_34_17_n_3392, mul_34_17_n_3393,
     mul_34_17_n_3394, mul_34_17_n_3395, mul_34_17_n_3396, mul_34_17_n_3397,
     mul_34_17_n_3398, mul_34_17_n_3399, mul_34_17_n_3400, mul_34_17_n_3401,
     mul_34_17_n_3402, mul_34_17_n_3403, mul_34_17_n_3404, mul_34_17_n_3405,
     mul_34_17_n_3406, mul_34_17_n_3407, mul_34_17_n_3408, mul_34_17_n_3409,
     mul_34_17_n_3410, mul_34_17_n_3411, mul_34_17_n_3412, mul_34_17_n_3413,
     mul_34_17_n_3414, mul_34_17_n_3415, mul_34_17_n_3416, mul_34_17_n_3417,
     mul_34_17_n_3418, mul_34_17_n_3419, mul_34_17_n_3420, mul_34_17_n_3421,
     mul_34_17_n_3422, mul_34_17_n_3423, mul_34_17_n_3424, mul_34_17_n_3425,
     mul_34_17_n_3426, mul_34_17_n_3427, mul_34_17_n_3428, mul_34_17_n_3429,
     mul_34_17_n_3430, mul_34_17_n_3431, mul_34_17_n_3432, mul_34_17_n_3433,
     mul_34_17_n_3434, mul_34_17_n_3435, mul_34_17_n_3436, mul_34_17_n_3437,
     mul_34_17_n_3438, mul_34_17_n_3439, mul_34_17_n_3440, mul_34_17_n_3441,
     mul_34_17_n_3442, mul_34_17_n_3443, mul_34_17_n_3444, mul_34_17_n_3445,
     mul_34_17_n_3446, mul_34_17_n_3447, mul_34_17_n_3448, mul_34_17_n_3449,
     mul_34_17_n_3450, mul_34_17_n_3451, mul_34_17_n_3452, mul_34_17_n_3453,
     mul_34_17_n_3454, mul_34_17_n_3455, mul_34_17_n_3456, mul_34_17_n_3457,
     mul_34_17_n_3458, mul_34_17_n_3459, mul_34_17_n_3460, mul_34_17_n_3461,
     mul_34_17_n_3462, mul_34_17_n_3463, mul_34_17_n_3464, mul_34_17_n_3465,
     mul_34_17_n_3466, mul_34_17_n_3467, mul_34_17_n_3468, mul_34_17_n_3469,
     mul_34_17_n_3470, mul_34_17_n_3471, mul_34_17_n_3472, mul_34_17_n_3473,
     mul_34_17_n_3474, mul_34_17_n_3475, mul_34_17_n_3476, mul_34_17_n_3477,
     mul_34_17_n_3478, mul_34_17_n_3479, mul_34_17_n_3480, mul_34_17_n_3481,
     mul_34_17_n_3482, mul_34_17_n_3483, mul_34_17_n_3484, mul_34_17_n_3485,
     mul_34_17_n_3486, mul_34_17_n_3487, mul_34_17_n_3488, mul_34_17_n_3489,
     mul_34_17_n_3490, mul_34_17_n_3491, mul_34_17_n_3492, mul_34_17_n_3493,
     mul_34_17_n_3494, mul_34_17_n_3495, mul_34_17_n_3496, mul_34_17_n_3497,
     mul_34_17_n_3498, mul_34_17_n_3499, mul_34_17_n_3500, mul_34_17_n_3501,
     mul_34_17_n_3502, mul_34_17_n_3503, mul_34_17_n_3504, mul_34_17_n_3505,
     mul_34_17_n_3506, mul_34_17_n_3507, mul_34_17_n_3508, mul_34_17_n_3509,
     mul_34_17_n_3510, mul_34_17_n_3511, mul_34_17_n_3512, mul_34_17_n_3513,
     mul_34_17_n_3514, mul_34_17_n_3515, mul_34_17_n_3516, mul_34_17_n_3517,
     mul_34_17_n_3518, mul_34_17_n_3519, mul_34_17_n_3520, mul_34_17_n_3521,
     mul_34_17_n_3522, mul_34_17_n_3523, mul_34_17_n_3524, mul_34_17_n_3525,
     mul_34_17_n_3526, mul_34_17_n_3527, mul_34_17_n_3528, mul_34_17_n_3529,
     mul_34_17_n_3530, mul_34_17_n_3531, mul_34_17_n_3532, mul_34_17_n_3533,
     mul_34_17_n_3534, mul_34_17_n_3535, mul_34_17_n_3536, mul_34_17_n_3537,
     mul_34_17_n_3538, mul_34_17_n_3539, mul_34_17_n_3540, mul_34_17_n_3541,
     mul_34_17_n_3542, mul_34_17_n_3543, mul_34_17_n_3544, mul_34_17_n_3545,
     mul_34_17_n_3546, mul_34_17_n_3547, mul_34_17_n_3548, mul_34_17_n_3549,
     mul_34_17_n_3550, mul_34_17_n_3551, mul_34_17_n_3552, mul_34_17_n_3553,
     mul_34_17_n_3554, mul_34_17_n_3555, mul_34_17_n_3556, mul_34_17_n_3557,
     mul_34_17_n_3558, mul_34_17_n_3559, mul_34_17_n_3560, mul_34_17_n_3561,
     mul_34_17_n_3562, mul_34_17_n_3563, mul_34_17_n_3564, mul_34_17_n_3565,
     mul_34_17_n_3566, mul_34_17_n_3567, mul_34_17_n_3568, mul_34_17_n_3569,
     mul_34_17_n_3570, mul_34_17_n_3571, mul_34_17_n_3572, mul_34_17_n_3573,
     mul_34_17_n_3574, mul_34_17_n_3575, mul_34_17_n_3576, mul_34_17_n_3577,
     mul_34_17_n_3578, mul_34_17_n_3579, mul_34_17_n_3580, mul_34_17_n_3581,
     mul_34_17_n_3582, mul_34_17_n_3583, mul_34_17_n_3584, mul_34_17_n_3585,
     mul_34_17_n_3586, mul_34_17_n_3587, mul_34_17_n_3588, mul_34_17_n_3589,
     mul_34_17_n_3590, mul_34_17_n_3591, mul_34_17_n_3592, mul_34_17_n_3593,
     mul_34_17_n_3594, mul_34_17_n_3595, mul_34_17_n_3596, mul_34_17_n_3597,
     mul_34_17_n_3598, mul_34_17_n_3599, mul_34_17_n_3600, mul_34_17_n_3601,
     mul_34_17_n_3602, mul_34_17_n_3603, mul_34_17_n_3604, mul_34_17_n_3605,
     mul_34_17_n_3606, mul_34_17_n_3607, mul_34_17_n_3608, mul_34_17_n_3609,
     mul_34_17_n_3610, mul_34_17_n_3611, mul_34_17_n_3612, mul_34_17_n_3613,
     mul_34_17_n_3614, mul_34_17_n_3615, mul_34_17_n_3616, mul_34_17_n_3617,
     mul_34_17_n_3618, mul_34_17_n_3619, mul_34_17_n_3620, mul_34_17_n_3621,
     mul_34_17_n_3622, mul_34_17_n_3623, mul_34_17_n_3624, mul_34_17_n_3625,
     mul_34_17_n_3626, mul_34_17_n_3627, mul_34_17_n_3628, mul_34_17_n_3629,
     mul_34_17_n_3630, mul_34_17_n_3631, mul_34_17_n_3632, mul_34_17_n_3633,
     mul_34_17_n_3634, mul_34_17_n_3635, mul_34_17_n_3636, mul_34_17_n_3637,
     mul_34_17_n_3638, mul_34_17_n_3639, mul_34_17_n_3640, mul_34_17_n_3641,
     mul_34_17_n_3642, mul_34_17_n_3643, mul_34_17_n_3644, mul_34_17_n_3645,
     mul_34_17_n_3646, mul_34_17_n_3647, mul_34_17_n_3648, mul_34_17_n_3649,
     mul_34_17_n_3650, mul_34_17_n_3651, mul_34_17_n_3652, mul_34_17_n_3653,
     mul_34_17_n_3654, mul_34_17_n_3655, mul_34_17_n_3656, mul_34_17_n_3657,
     mul_34_17_n_3658, mul_34_17_n_3659, mul_34_17_n_3660, mul_34_17_n_3661,
     mul_34_17_n_3662, mul_34_17_n_3663, mul_34_17_n_3664, mul_34_17_n_3665,
     mul_34_17_n_3666, mul_34_17_n_3667, mul_34_17_n_3668, mul_34_17_n_3669,
     mul_34_17_n_3670, mul_34_17_n_3671, mul_34_17_n_3672, mul_34_17_n_3673,
     mul_34_17_n_3674, mul_34_17_n_3675, mul_34_17_n_3676, mul_34_17_n_3677,
     mul_34_17_n_3678, mul_34_17_n_3679, mul_34_17_n_3680, mul_34_17_n_3681,
     mul_34_17_n_3682, mul_34_17_n_3683, mul_34_17_n_3684, mul_34_17_n_3685,
     mul_34_17_n_3686, mul_34_17_n_3687, mul_34_17_n_3688, mul_34_17_n_3689,
     mul_34_17_n_3690, mul_34_17_n_3691, mul_34_17_n_3692, mul_34_17_n_3693,
     mul_34_17_n_3694, mul_34_17_n_3695, mul_34_17_n_3696, mul_34_17_n_3697,
     mul_34_17_n_3698, mul_34_17_n_3699, mul_34_17_n_3700, mul_34_17_n_3701,
     mul_34_17_n_3702, mul_34_17_n_3703, mul_34_17_n_3704, mul_34_17_n_3705,
     mul_34_17_n_3706, mul_34_17_n_3707, mul_34_17_n_3708, mul_34_17_n_3709,
     mul_34_17_n_3710, mul_34_17_n_3711, mul_34_17_n_3712, mul_34_17_n_3713,
     mul_34_17_n_3714, mul_34_17_n_3715, mul_34_17_n_3716, mul_34_17_n_3717,
     mul_34_17_n_3718, mul_34_17_n_3719, mul_34_17_n_3720, mul_34_17_n_3721,
     mul_34_17_n_3722, mul_34_17_n_3723, mul_34_17_n_3724, mul_34_17_n_3725,
     mul_34_17_n_3726, mul_34_17_n_3727, mul_34_17_n_3728, mul_34_17_n_3729,
     mul_34_17_n_3730, mul_34_17_n_3731, mul_34_17_n_3732, mul_34_17_n_3733,
     mul_34_17_n_3734, mul_34_17_n_3735, mul_34_17_n_3736, mul_34_17_n_3737,
     mul_34_17_n_3738, mul_34_17_n_3739, mul_34_17_n_3740, mul_34_17_n_3741,
     mul_34_17_n_3742, mul_34_17_n_3743, mul_34_17_n_3744, mul_34_17_n_3745,
     mul_34_17_n_3746, mul_34_17_n_3747, mul_34_17_n_3748, mul_34_17_n_3749,
     mul_34_17_n_3750, mul_34_17_n_3751, mul_34_17_n_3752, mul_34_17_n_3753,
     mul_34_17_n_3754, mul_34_17_n_3755, mul_34_17_n_3756, mul_34_17_n_3757,
     mul_34_17_n_3758, mul_34_17_n_3759, mul_34_17_n_3760, mul_34_17_n_3761,
     mul_34_17_n_3762, mul_34_17_n_3763, mul_34_17_n_3764, mul_34_17_n_3765,
     mul_34_17_n_3766, mul_34_17_n_3767, mul_34_17_n_3768, mul_34_17_n_3769,
     mul_34_17_n_3770, mul_34_17_n_3771, mul_34_17_n_3772, mul_34_17_n_3773,
     mul_34_17_n_3774, mul_34_17_n_3775, mul_34_17_n_3776, mul_34_17_n_3777,
     mul_34_17_n_3778, mul_34_17_n_3779, mul_34_17_n_3780, mul_34_17_n_3781,
     mul_34_17_n_3782, mul_34_17_n_3783, mul_34_17_n_3784, mul_34_17_n_3785,
     mul_34_17_n_3786, mul_34_17_n_3787, mul_34_17_n_3788, mul_34_17_n_3789,
     mul_34_17_n_3790, mul_34_17_n_3791, mul_34_17_n_3792, mul_34_17_n_3793,
     mul_34_17_n_3794, mul_34_17_n_3795, mul_34_17_n_3796, mul_34_17_n_3797,
     mul_34_17_n_3798, mul_34_17_n_3799, mul_34_17_n_3800, mul_34_17_n_3801,
     mul_34_17_n_3802, mul_34_17_n_3803, mul_34_17_n_3804, mul_34_17_n_3805,
     mul_34_17_n_3806, mul_34_17_n_3807, mul_34_17_n_3808, mul_34_17_n_3809,
     mul_34_17_n_3810, mul_34_17_n_3811, mul_34_17_n_3812, mul_34_17_n_3813,
     mul_34_17_n_3814, mul_34_17_n_3815, mul_34_17_n_3816, mul_34_17_n_3817,
     mul_34_17_n_3818, mul_34_17_n_3819, mul_34_17_n_3820, mul_34_17_n_3821,
     mul_34_17_n_3822, mul_34_17_n_3823, mul_34_17_n_3824, mul_34_17_n_3825,
     mul_34_17_n_3826, mul_34_17_n_3827, mul_34_17_n_3828, mul_34_17_n_3829,
     mul_34_17_n_3830, mul_34_17_n_3831, mul_34_17_n_3832, mul_34_17_n_3833,
     mul_34_17_n_3834, mul_34_17_n_3835, mul_34_17_n_3836, mul_34_17_n_3837,
     mul_34_17_n_3838, mul_34_17_n_3839, mul_34_17_n_3840, mul_34_17_n_3841,
     mul_34_17_n_3842, mul_34_17_n_3843, mul_34_17_n_3844, mul_34_17_n_3845,
     mul_34_17_n_3846, mul_34_17_n_3847, mul_34_17_n_3848, mul_34_17_n_3849,
     mul_34_17_n_3850, mul_34_17_n_3851, mul_34_17_n_3852, mul_34_17_n_3853,
     mul_34_17_n_3854, mul_34_17_n_3855, mul_34_17_n_3856, mul_34_17_n_3857,
     mul_34_17_n_3858, mul_34_17_n_3859, mul_34_17_n_3860, mul_34_17_n_3861,
     mul_34_17_n_3862, mul_34_17_n_3863, mul_34_17_n_3864, mul_34_17_n_3865,
     mul_34_17_n_3866, mul_34_17_n_3867, mul_34_17_n_3868, mul_34_17_n_3869,
     mul_34_17_n_3870, mul_34_17_n_3871, mul_34_17_n_3872, mul_34_17_n_3873,
     mul_34_17_n_3874, mul_34_17_n_3875, mul_34_17_n_3876, mul_34_17_n_3877,
     mul_34_17_n_3878, mul_34_17_n_3879, mul_34_17_n_3880, mul_34_17_n_3881,
     mul_34_17_n_3882, mul_34_17_n_3883, mul_34_17_n_3884, mul_34_17_n_3885,
     mul_34_17_n_3886, mul_34_17_n_3887, mul_34_17_n_3888, mul_34_17_n_3889,
     mul_34_17_n_3890, mul_34_17_n_3891, mul_34_17_n_3892, mul_34_17_n_3893,
     mul_34_17_n_3894, mul_34_17_n_3895, mul_34_17_n_3896, mul_34_17_n_3897,
     mul_34_17_n_3898, mul_34_17_n_3899, mul_34_17_n_3900, mul_34_17_n_3901,
     mul_34_17_n_3902, mul_34_17_n_3903, mul_34_17_n_3904, mul_34_17_n_3905,
     mul_34_17_n_3906, mul_34_17_n_3907, mul_34_17_n_3908, mul_34_17_n_3909,
     mul_34_17_n_3910, mul_34_17_n_3911, mul_34_17_n_3912, mul_34_17_n_3913,
     mul_34_17_n_3914, mul_34_17_n_3915, mul_34_17_n_3916, mul_34_17_n_3917,
     mul_34_17_n_3918, mul_34_17_n_3919, mul_34_17_n_3920, mul_34_17_n_3921,
     mul_34_17_n_3922, mul_34_17_n_3923, mul_34_17_n_3924, mul_34_17_n_3925,
     mul_34_17_n_3926, mul_34_17_n_3927, mul_34_17_n_3928, mul_34_17_n_3929,
     mul_34_17_n_3930, mul_34_17_n_3931, mul_34_17_n_3932, mul_34_17_n_3933,
     mul_34_17_n_3934, mul_34_17_n_3935, mul_34_17_n_3936, mul_34_17_n_3937,
     mul_34_17_n_3938, mul_34_17_n_3939, mul_34_17_n_3940, mul_34_17_n_3941,
     mul_34_17_n_3942, mul_34_17_n_3943, mul_34_17_n_3944, mul_34_17_n_3945,
     mul_34_17_n_3946, mul_34_17_n_3947, mul_34_17_n_3948, mul_34_17_n_3949,
     mul_34_17_n_3950, mul_34_17_n_3951, mul_34_17_n_3952, mul_34_17_n_3953,
     mul_34_17_n_3954, mul_34_17_n_3955, mul_34_17_n_3956, mul_34_17_n_3957,
     mul_34_17_n_3958, mul_34_17_n_3959, mul_34_17_n_3960, mul_34_17_n_3961,
     mul_34_17_n_3962, mul_34_17_n_3963, mul_34_17_n_3964, mul_34_17_n_3965,
     mul_34_17_n_3966, mul_34_17_n_3967, mul_34_17_n_3968, mul_34_17_n_3969,
     mul_34_17_n_3970, mul_34_17_n_3971, mul_34_17_n_3972, mul_34_17_n_3973,
     mul_34_17_n_3974, mul_34_17_n_3975, mul_34_17_n_3976, mul_34_17_n_3977,
     mul_34_17_n_3978, mul_34_17_n_3979, mul_34_17_n_3980, mul_34_17_n_3981,
     mul_34_17_n_3982, mul_34_17_n_3983, mul_34_17_n_3984, mul_34_17_n_3985,
     mul_34_17_n_3986, mul_34_17_n_3987, mul_34_17_n_3988, mul_34_17_n_3989,
     mul_34_17_n_3990, mul_34_17_n_3991, mul_34_17_n_3992, mul_34_17_n_3993,
     mul_34_17_n_3994, mul_34_17_n_3995, mul_34_17_n_3996, mul_34_17_n_3997,
     mul_34_17_n_3998, mul_34_17_n_3999, mul_34_17_n_4000, mul_34_17_n_4001,
     mul_34_17_n_4002, mul_34_17_n_4003, mul_34_17_n_4004, mul_34_17_n_4005,
     mul_34_17_n_4006, mul_34_17_n_4007, mul_34_17_n_4008, mul_34_17_n_4009,
     mul_34_17_n_4010, mul_34_17_n_4011, mul_34_17_n_4012, mul_34_17_n_4013,
     mul_34_17_n_4014, mul_34_17_n_4015, mul_34_17_n_4016, mul_34_17_n_4017,
     mul_34_17_n_4018, mul_34_17_n_4019, mul_34_17_n_4020, mul_34_17_n_4021,
     mul_34_17_n_4022, mul_34_17_n_4023, mul_34_17_n_4024, mul_34_17_n_4025,
     mul_34_17_n_4026, mul_34_17_n_4027, mul_34_17_n_4028, mul_34_17_n_4029,
     mul_34_17_n_4030, mul_34_17_n_4031, mul_34_17_n_4032, mul_34_17_n_4033,
     mul_34_17_n_4034, mul_34_17_n_4035, mul_34_17_n_4036, mul_34_17_n_4037,
     mul_34_17_n_4038, mul_34_17_n_4039, mul_34_17_n_4040, mul_34_17_n_4041,
     mul_34_17_n_4042, mul_34_17_n_4043, mul_34_17_n_4044, mul_34_17_n_4045,
     mul_34_17_n_4046, mul_34_17_n_4047, mul_34_17_n_4048, mul_34_17_n_4049,
     mul_34_17_n_4050, mul_34_17_n_4051, mul_34_17_n_4052, mul_34_17_n_4053,
     mul_34_17_n_4054, mul_34_17_n_4055, mul_34_17_n_4056, mul_34_17_n_4057,
     mul_34_17_n_4058, mul_34_17_n_4059, mul_34_17_n_4060, mul_34_17_n_4061,
     mul_34_17_n_4062, mul_34_17_n_4063, mul_34_17_n_4064, mul_34_17_n_4065,
     mul_34_17_n_4066, mul_34_17_n_4067, mul_34_17_n_4068, mul_34_17_n_4069,
     mul_34_17_n_4070, mul_34_17_n_4071, mul_34_17_n_4072, mul_34_17_n_4073,
     mul_34_17_n_4074, mul_34_17_n_4075, mul_34_17_n_4076, mul_34_17_n_4077,
     mul_34_17_n_4078, mul_34_17_n_4079, mul_34_17_n_4080, mul_34_17_n_4081,
     mul_34_17_n_4082, mul_34_17_n_4083, mul_34_17_n_4084, mul_34_17_n_4085,
     mul_34_17_n_4086, mul_34_17_n_4087, mul_34_17_n_4088, mul_34_17_n_4089,
     mul_34_17_n_4090, mul_34_17_n_4091, mul_34_17_n_4092, mul_34_17_n_4093,
     mul_34_17_n_4094, mul_34_17_n_4095, mul_34_17_n_4096, mul_34_17_n_4097,
     mul_34_17_n_4098, mul_34_17_n_4099, mul_34_17_n_4100, mul_34_17_n_4101,
     mul_34_17_n_4102, mul_34_17_n_4103, mul_34_17_n_4104, mul_34_17_n_4105,
     mul_34_17_n_4106, mul_34_17_n_4107, mul_34_17_n_4108, mul_34_17_n_4109,
     mul_34_17_n_4110, mul_34_17_n_4111, mul_34_17_n_4112, mul_34_17_n_4113,
     mul_34_17_n_4114, mul_34_17_n_4115, mul_34_17_n_4116, mul_34_17_n_4117,
     mul_34_17_n_4118, mul_34_17_n_4119, mul_34_17_n_4120, mul_34_17_n_4121,
     mul_34_17_n_4122, mul_34_17_n_4123, mul_34_17_n_4124, mul_34_17_n_4125,
     mul_34_17_n_4126, mul_34_17_n_4127, mul_34_17_n_4128, mul_34_17_n_4129,
     mul_34_17_n_4130, mul_34_17_n_4131, mul_34_17_n_4132, mul_34_17_n_4133,
     mul_34_17_n_4134, mul_34_17_n_4135, mul_34_17_n_4136, mul_34_17_n_4137,
     mul_34_17_n_4138, mul_34_17_n_4139, mul_34_17_n_4140, mul_34_17_n_4141,
     mul_34_17_n_4142, mul_34_17_n_4143, mul_34_17_n_4144, mul_34_17_n_4145,
     mul_34_17_n_4146, mul_34_17_n_4147, mul_34_17_n_4148, mul_34_17_n_4149,
     mul_34_17_n_4150, mul_34_17_n_4151, mul_34_17_n_4152, mul_34_17_n_4153,
     mul_34_17_n_4154, mul_34_17_n_4155, mul_34_17_n_4156, mul_34_17_n_4157,
     mul_34_17_n_4158, mul_34_17_n_4159, mul_34_17_n_4160, mul_34_17_n_4161,
     mul_34_17_n_4162, mul_34_17_n_4163, mul_34_17_n_4164, mul_34_17_n_4165,
     mul_34_17_n_4166, mul_34_17_n_4167, mul_34_17_n_4168, mul_34_17_n_4169,
     mul_34_17_n_4170, mul_34_17_n_4171, mul_34_17_n_4172, mul_34_17_n_4173,
     mul_34_17_n_4174, mul_34_17_n_4175, mul_34_17_n_4176, mul_34_17_n_4177,
     mul_34_17_n_4178, mul_34_17_n_4179, mul_34_17_n_4180, mul_34_17_n_4181,
     mul_34_17_n_4182, mul_34_17_n_4183, mul_34_17_n_4184, mul_34_17_n_4185,
     mul_34_17_n_4186, mul_34_17_n_4187, mul_34_17_n_4188, mul_34_17_n_4189,
     mul_34_17_n_4190, mul_34_17_n_4191, mul_34_17_n_4192, mul_34_17_n_4193,
     mul_34_17_n_4194, mul_34_17_n_4195, mul_34_17_n_4196, mul_34_17_n_4197,
     mul_34_17_n_4198, mul_34_17_n_4199, mul_34_17_n_4200, mul_34_17_n_4201,
     mul_34_17_n_4202, mul_34_17_n_4203, mul_34_17_n_4204, mul_34_17_n_4205,
     mul_34_17_n_4206, mul_34_17_n_4207, mul_34_17_n_4208, mul_34_17_n_4209,
     mul_34_17_n_4210, mul_34_17_n_4211, mul_34_17_n_4212, mul_34_17_n_4213,
     mul_34_17_n_4214, mul_34_17_n_4215, mul_34_17_n_4216, mul_34_17_n_4217,
     mul_34_17_n_4218, mul_34_17_n_4219, mul_34_17_n_4220, mul_34_17_n_4221,
     mul_34_17_n_4222, mul_34_17_n_4223, mul_34_17_n_4224, mul_34_17_n_4225,
     mul_34_17_n_4226, mul_34_17_n_4227, mul_34_17_n_4228, mul_34_17_n_4229,
     mul_34_17_n_4230, mul_34_17_n_4231, mul_34_17_n_4232, mul_34_17_n_4233,
     mul_34_17_n_4234, mul_34_17_n_4235, mul_34_17_n_4236, mul_34_17_n_4237,
     mul_34_17_n_4238, mul_34_17_n_4239, mul_34_17_n_4240, mul_34_17_n_4241,
     mul_34_17_n_4242, mul_34_17_n_4243, mul_34_17_n_4244, mul_34_17_n_4245,
     mul_34_17_n_4246, mul_34_17_n_4247, mul_34_17_n_4248, mul_34_17_n_4249,
     mul_34_17_n_4250, mul_34_17_n_4251, mul_34_17_n_4252, mul_34_17_n_4253,
     mul_34_17_n_4254, mul_34_17_n_4255, mul_34_17_n_4256, mul_34_17_n_4257,
     mul_34_17_n_4258, mul_34_17_n_4259, mul_34_17_n_4260, mul_34_17_n_4261,
     mul_34_17_n_4262, mul_34_17_n_4263, mul_34_17_n_4264, mul_34_17_n_4265,
     mul_34_17_n_4266, mul_34_17_n_4267, mul_34_17_n_4268, mul_34_17_n_4269,
     mul_34_17_n_4270, mul_34_17_n_4271, mul_34_17_n_4272, mul_34_17_n_4273,
     mul_34_17_n_4274, mul_34_17_n_4275, mul_34_17_n_4276, mul_34_17_n_4277,
     mul_34_17_n_4278, mul_34_17_n_4279, mul_34_17_n_4280, mul_34_17_n_4281,
     mul_34_17_n_4282, mul_34_17_n_4283, mul_34_17_n_4284, mul_34_17_n_4285,
     mul_34_17_n_4286, mul_34_17_n_4287, mul_34_17_n_4288, mul_34_17_n_4289,
     mul_34_17_n_4290, mul_34_17_n_4291, mul_34_17_n_4292, mul_34_17_n_4293,
     mul_34_17_n_4294, mul_34_17_n_4295, mul_34_17_n_4296, mul_34_17_n_4297,
     mul_34_17_n_4298, mul_34_17_n_4299, mul_34_17_n_4300, mul_34_17_n_4301,
     mul_34_17_n_4302, mul_34_17_n_4303, mul_34_17_n_4304, mul_34_17_n_4305,
     mul_34_17_n_4306, mul_34_17_n_4307, mul_34_17_n_4308, mul_34_17_n_4309,
     mul_34_17_n_4310, mul_34_17_n_4311, mul_34_17_n_4312, mul_34_17_n_4313,
     mul_34_17_n_4314, mul_34_17_n_4315, mul_34_17_n_4316, mul_34_17_n_4317,
     mul_34_17_n_4318, mul_34_17_n_4319, mul_34_17_n_4320, mul_34_17_n_4321,
     mul_34_17_n_4322, mul_34_17_n_4323, mul_34_17_n_4324, mul_34_17_n_4325,
     mul_34_17_n_4326, mul_34_17_n_4327, mul_34_17_n_4328, mul_34_17_n_4329,
     mul_34_17_n_4330, mul_34_17_n_4331, mul_34_17_n_4332, mul_34_17_n_4333,
     mul_34_17_n_4334, mul_34_17_n_4335, mul_34_17_n_4336, mul_34_17_n_4337,
     mul_34_17_n_4338, mul_34_17_n_4339, mul_34_17_n_4340, mul_34_17_n_4341,
     mul_34_17_n_4342, mul_34_17_n_4343, mul_34_17_n_4344, mul_34_17_n_4345,
     mul_34_17_n_4346, mul_34_17_n_4347, mul_34_17_n_4348, mul_34_17_n_4349,
     mul_34_17_n_4350, mul_34_17_n_4351, mul_34_17_n_4352, mul_34_17_n_4353,
     mul_34_17_n_4354, mul_34_17_n_4355, mul_34_17_n_4356, mul_34_17_n_4357,
     mul_34_17_n_4358, mul_34_17_n_4359, mul_34_17_n_4360, mul_34_17_n_4361,
     mul_34_17_n_4362, mul_34_17_n_4363, mul_34_17_n_4364, mul_34_17_n_4365,
     mul_34_17_n_4366, mul_34_17_n_4367, mul_34_17_n_4368, mul_34_17_n_4369,
     mul_34_17_n_4370, mul_34_17_n_4371, mul_34_17_n_4372, mul_34_17_n_4373,
     mul_34_17_n_4374, mul_34_17_n_4375, mul_34_17_n_4376, mul_34_17_n_4377,
     mul_34_17_n_4378, mul_34_17_n_4379, mul_34_17_n_4380, mul_34_17_n_4381,
     mul_34_17_n_4382, mul_34_17_n_4383, mul_34_17_n_4384, mul_34_17_n_4385,
     mul_34_17_n_4386, mul_34_17_n_4387, mul_34_17_n_4388, mul_34_17_n_4389,
     mul_34_17_n_4390, mul_34_17_n_4391, mul_34_17_n_4392, mul_34_17_n_4393,
     mul_34_17_n_4394, mul_34_17_n_4395, mul_34_17_n_4396, mul_34_17_n_4397,
     mul_34_17_n_4398, mul_34_17_n_4399, mul_34_17_n_4400, mul_34_17_n_4401,
     mul_34_17_n_4402, mul_34_17_n_4403, mul_34_17_n_4404, mul_34_17_n_4405,
     mul_34_17_n_4406, mul_34_17_n_4407, mul_34_17_n_4408, mul_34_17_n_4409,
     mul_34_17_n_4410, mul_34_17_n_4411, mul_34_17_n_4412, mul_34_17_n_4413,
     mul_34_17_n_4414, mul_34_17_n_4415, mul_34_17_n_4416, mul_34_17_n_4417,
     mul_34_17_n_4418, mul_34_17_n_4419, mul_34_17_n_4420, mul_34_17_n_4421,
     mul_34_17_n_4422, mul_34_17_n_4423, mul_34_17_n_4424, mul_34_17_n_4425,
     mul_34_17_n_4426, mul_34_17_n_4427, mul_34_17_n_4428, mul_34_17_n_4429,
     mul_34_17_n_4430, mul_34_17_n_4431, mul_34_17_n_4432, mul_34_17_n_4433,
     mul_34_17_n_4434, mul_34_17_n_4435, mul_34_17_n_4436, mul_34_17_n_4437,
     mul_34_17_n_4438, mul_34_17_n_4439, mul_34_17_n_4440, mul_34_17_n_4441,
     mul_34_17_n_4442, mul_34_17_n_4443, mul_34_17_n_4444, mul_34_17_n_4445,
     mul_34_17_n_4446, mul_34_17_n_4447, mul_34_17_n_4448, mul_34_17_n_4449,
     mul_34_17_n_4450, mul_34_17_n_4451, mul_34_17_n_4452, mul_34_17_n_4453,
     mul_34_17_n_4454, mul_34_17_n_4455, mul_34_17_n_4456, mul_34_17_n_4457,
     mul_34_17_n_4458, mul_34_17_n_4459, mul_34_17_n_4460, mul_34_17_n_4461,
     mul_34_17_n_4462, mul_34_17_n_4463, mul_34_17_n_4464, mul_34_17_n_4465,
     mul_34_17_n_4466, mul_34_17_n_4467, mul_34_17_n_4468, mul_34_17_n_4469,
     mul_34_17_n_4470, mul_34_17_n_4471, mul_34_17_n_4472, mul_34_17_n_4473,
     mul_34_17_n_4474, mul_34_17_n_4475, mul_34_17_n_4476, mul_34_17_n_4477,
     mul_34_17_n_4478, mul_34_17_n_4479, mul_34_17_n_4480, mul_34_17_n_4481,
     mul_34_17_n_4482, mul_34_17_n_4483, mul_34_17_n_4484, mul_34_17_n_4485,
     mul_34_17_n_4486, mul_34_17_n_4487, mul_34_17_n_4488, mul_34_17_n_4489,
     mul_34_17_n_4490, mul_34_17_n_4491, mul_34_17_n_4492, mul_34_17_n_4493,
     mul_34_17_n_4494, mul_34_17_n_4495, mul_34_17_n_4496, mul_34_17_n_4497,
     mul_34_17_n_4498, mul_34_17_n_4499, mul_34_17_n_4500, mul_34_17_n_4501,
     mul_34_17_n_4502, mul_34_17_n_4503, mul_34_17_n_4504, mul_34_17_n_4505,
     mul_34_17_n_4506, mul_34_17_n_4507, mul_34_17_n_4508, mul_34_17_n_4509,
     mul_34_17_n_4510, mul_34_17_n_4511, mul_34_17_n_4512, mul_34_17_n_4513,
     mul_34_17_n_4514, mul_34_17_n_4515, mul_34_17_n_4516, mul_34_17_n_4517,
     mul_34_17_n_4518, mul_34_17_n_4519, mul_34_17_n_4520, mul_34_17_n_4521,
     mul_34_17_n_4522, mul_34_17_n_4523, mul_34_17_n_4524, mul_34_17_n_4525,
     mul_34_17_n_4526, mul_34_17_n_4527, mul_34_17_n_4528, mul_34_17_n_4529,
     mul_34_17_n_4530, mul_34_17_n_4531, mul_34_17_n_4532, mul_34_17_n_4533,
     mul_34_17_n_4534, mul_34_17_n_4535, mul_34_17_n_4536, mul_34_17_n_4537,
     mul_34_17_n_4538, mul_34_17_n_4539, mul_34_17_n_4540, mul_34_17_n_4541,
     mul_34_17_n_4542, mul_34_17_n_4543, mul_34_17_n_4544, mul_34_17_n_4545,
     mul_34_17_n_4546, mul_34_17_n_4547, mul_34_17_n_4548, mul_34_17_n_4549,
     mul_34_17_n_4550, mul_34_17_n_4551, mul_34_17_n_4552, mul_34_17_n_4553,
     mul_34_17_n_4554, mul_34_17_n_4555, mul_34_17_n_4556, mul_34_17_n_4557,
     mul_34_17_n_4558, mul_34_17_n_4559, mul_34_17_n_4560, mul_34_17_n_4561,
     mul_34_17_n_4562, mul_34_17_n_4563, mul_34_17_n_4564, mul_34_17_n_4565,
     mul_34_17_n_4566, mul_34_17_n_4567, mul_34_17_n_4568, mul_34_17_n_4569,
     mul_34_17_n_4570, mul_34_17_n_4571, mul_34_17_n_4572, mul_34_17_n_4573,
     mul_34_17_n_4574, mul_34_17_n_4575, mul_34_17_n_4576, mul_34_17_n_4577,
     mul_34_17_n_4578, mul_34_17_n_4579, mul_34_17_n_4580, mul_34_17_n_4581,
     mul_34_17_n_4582, mul_34_17_n_4583, mul_34_17_n_4584, mul_34_17_n_4585,
     mul_34_17_n_4586, mul_34_17_n_4587, mul_34_17_n_4588, mul_34_17_n_4589,
     mul_34_17_n_4590, mul_34_17_n_4591, mul_34_17_n_4592, mul_34_17_n_4593,
     mul_34_17_n_4594, mul_34_17_n_4595, mul_34_17_n_4596, mul_34_17_n_4597,
     mul_34_17_n_4598, mul_34_17_n_4599, mul_34_17_n_4600, mul_34_17_n_4601,
     mul_34_17_n_4602, mul_34_17_n_4603, mul_34_17_n_4604, mul_34_17_n_4605,
     mul_34_17_n_4606, mul_34_17_n_4607, mul_34_17_n_4608, mul_34_17_n_4609,
     mul_34_17_n_4610, mul_34_17_n_4611, mul_34_17_n_4612, mul_34_17_n_4613,
     mul_34_17_n_4614, mul_34_17_n_4615, mul_34_17_n_4616, mul_34_17_n_4617,
     mul_34_17_n_4618, mul_34_17_n_4619, mul_34_17_n_4620, mul_34_17_n_4621,
     mul_34_17_n_4622, mul_34_17_n_4623, mul_34_17_n_4624, mul_34_17_n_4625,
     mul_34_17_n_4626, mul_34_17_n_4627, mul_34_17_n_4628, mul_34_17_n_4629,
     mul_34_17_n_4630, mul_34_17_n_4631, mul_34_17_n_4632, mul_34_17_n_4633,
     mul_34_17_n_4634, mul_34_17_n_4635, mul_34_17_n_4636, mul_34_17_n_4637,
     mul_34_17_n_4638, mul_34_17_n_4639, mul_34_17_n_4640, mul_34_17_n_4641,
     mul_34_17_n_4642, mul_34_17_n_4643, mul_34_17_n_4644, mul_34_17_n_4645,
     mul_34_17_n_4646, mul_34_17_n_4647, mul_34_17_n_4648, mul_34_17_n_4649,
     mul_34_17_n_4650, mul_34_17_n_4651, mul_34_17_n_4652, mul_34_17_n_4653,
     mul_34_17_n_4654, mul_34_17_n_4655, mul_34_17_n_4656, mul_34_17_n_4657,
     mul_34_17_n_4658, mul_34_17_n_4659, mul_34_17_n_4660, mul_34_17_n_4661,
     mul_34_17_n_4662, mul_34_17_n_4663, mul_34_17_n_4664, mul_34_17_n_4665,
     mul_34_17_n_4666, mul_34_17_n_4667, mul_34_17_n_4668, mul_34_17_n_4669,
     mul_34_17_n_4670, mul_34_17_n_4671, mul_34_17_n_4672, mul_34_17_n_4673,
     mul_34_17_n_4674, mul_34_17_n_4675, mul_34_17_n_4676, mul_34_17_n_4677,
     mul_34_17_n_4678, mul_34_17_n_4679, mul_34_17_n_4680, mul_34_17_n_4681,
     mul_34_17_n_4682, mul_34_17_n_4683, mul_34_17_n_4684, mul_34_17_n_4685,
     mul_34_17_n_4686, mul_34_17_n_4687, mul_34_17_n_4688, mul_34_17_n_4689,
     mul_34_17_n_4690, mul_34_17_n_4691, mul_34_17_n_4692, mul_34_17_n_4693,
     mul_34_17_n_4694, mul_34_17_n_4695, mul_34_17_n_4696, mul_34_17_n_4697,
     mul_34_17_n_4698, mul_34_17_n_4699, mul_34_17_n_4700, mul_34_17_n_4701,
     mul_34_17_n_4702, mul_34_17_n_4703, mul_34_17_n_4704, mul_34_17_n_4705,
     mul_34_17_n_4706, mul_34_17_n_4707, mul_34_17_n_4708, mul_34_17_n_4709,
     mul_34_17_n_4710, mul_34_17_n_4711, mul_34_17_n_4712, mul_34_17_n_4713,
     mul_34_17_n_4714, mul_34_17_n_4715, mul_34_17_n_4716, mul_34_17_n_4717,
     mul_34_17_n_4718, mul_34_17_n_4719, mul_34_17_n_4720, mul_34_17_n_4721,
     mul_34_17_n_4722, mul_34_17_n_4723, mul_34_17_n_4724, mul_34_17_n_4725,
     mul_34_17_n_4726, mul_34_17_n_4727, mul_34_17_n_4728, mul_34_17_n_4729,
     mul_34_17_n_4730, mul_34_17_n_4731, mul_34_17_n_4732, mul_34_17_n_4733,
     mul_34_17_n_4734, mul_34_17_n_4735, mul_34_17_n_4736, mul_34_17_n_4737,
     mul_34_17_n_4738, mul_34_17_n_4739, mul_34_17_n_4740, mul_34_17_n_4741,
     mul_34_17_n_4742, mul_34_17_n_4743, mul_34_17_n_4744, mul_34_17_n_4745,
     mul_34_17_n_4746, mul_34_17_n_4747, mul_34_17_n_4748, mul_34_17_n_4749,
     mul_34_17_n_4750, mul_34_17_n_4751, mul_34_17_n_4752, mul_34_17_n_4753,
     mul_34_17_n_4754, mul_34_17_n_4755, mul_34_17_n_4756, mul_34_17_n_4757,
     mul_34_17_n_4758, mul_34_17_n_4759, mul_34_17_n_4760, mul_34_17_n_4761,
     mul_34_17_n_4762, mul_34_17_n_4763, mul_34_17_n_4764, mul_34_17_n_4765,
     mul_34_17_n_4766, mul_34_17_n_4767, mul_34_17_n_4768, mul_34_17_n_4769,
     mul_34_17_n_4770, mul_34_17_n_4771, mul_34_17_n_4772, mul_34_17_n_4773,
     mul_34_17_n_4774, mul_34_17_n_4775, mul_34_17_n_4776, mul_34_17_n_4777,
     mul_34_17_n_4778, mul_34_17_n_4779, mul_34_17_n_4780, mul_34_17_n_4781,
     mul_34_17_n_4782, mul_34_17_n_4783, mul_34_17_n_4784, mul_34_17_n_4785,
     mul_34_17_n_4786, mul_34_17_n_4787, mul_34_17_n_4788, mul_34_17_n_4789,
     mul_34_17_n_4790, mul_34_17_n_4791, mul_34_17_n_4792, mul_34_17_n_4793,
     mul_34_17_n_4794, mul_34_17_n_4795, mul_34_17_n_4796, mul_34_17_n_4797,
     mul_34_17_n_4798, mul_34_17_n_4799, mul_34_17_n_4800, mul_34_17_n_4801,
     mul_34_17_n_4802, mul_34_17_n_4803, mul_34_17_n_4804, mul_34_17_n_4805,
     mul_34_17_n_4806, mul_34_17_n_4807, mul_34_17_n_4808, mul_34_17_n_4809,
     mul_34_17_n_4810, mul_34_17_n_4811, mul_34_17_n_4812, mul_34_17_n_4813,
     mul_34_17_n_4814, mul_34_17_n_4815, mul_34_17_n_4816, mul_34_17_n_4817,
     mul_34_17_n_4818, mul_34_17_n_4819, mul_34_17_n_4820, mul_34_17_n_4821,
     mul_34_17_n_4822, mul_34_17_n_4823, mul_34_17_n_4824, mul_34_17_n_4825,
     mul_34_17_n_4826, mul_34_17_n_4827, mul_34_17_n_4828, mul_34_17_n_4829,
     mul_34_17_n_4830, mul_34_17_n_4831, mul_34_17_n_4832, mul_34_17_n_4833,
     mul_34_17_n_4834, mul_34_17_n_4835, mul_34_17_n_4836, mul_34_17_n_4837,
     mul_34_17_n_4838, mul_34_17_n_4839, mul_34_17_n_4840, mul_34_17_n_4841,
     mul_34_17_n_4842, mul_34_17_n_4843, mul_34_17_n_4844, mul_34_17_n_4845,
     mul_34_17_n_4846, mul_34_17_n_4847, mul_34_17_n_4848, mul_34_17_n_4849,
     mul_34_17_n_4850, mul_34_17_n_4851, mul_34_17_n_4852, mul_34_17_n_4853,
     mul_34_17_n_4854, mul_34_17_n_4855, mul_34_17_n_4856, mul_34_17_n_4857,
     mul_34_17_n_4858, mul_34_17_n_4859, mul_34_17_n_4860, mul_34_17_n_4861,
     mul_34_17_n_4862, mul_34_17_n_4863, mul_34_17_n_4864, mul_34_17_n_4865,
     mul_34_17_n_4866, mul_34_17_n_4867, mul_34_17_n_4868, mul_34_17_n_4869,
     mul_34_17_n_4870, mul_34_17_n_4871, mul_34_17_n_4872, mul_34_17_n_4873,
     mul_34_17_n_4874, mul_34_17_n_4875, mul_34_17_n_4876, mul_34_17_n_4877,
     mul_34_17_n_4878, mul_34_17_n_4879, mul_34_17_n_4880, mul_34_17_n_4881,
     mul_34_17_n_4882, mul_34_17_n_4883, mul_34_17_n_4884, mul_34_17_n_4885,
     mul_34_17_n_4886, mul_34_17_n_4887, mul_34_17_n_4888, mul_34_17_n_4889,
     mul_34_17_n_4890, mul_34_17_n_4891, mul_34_17_n_4892, mul_34_17_n_4893,
     mul_34_17_n_4894, mul_34_17_n_4895, mul_34_17_n_4896, mul_34_17_n_4897,
     mul_34_17_n_4898, mul_34_17_n_4899, mul_34_17_n_4900, mul_34_17_n_4901,
     mul_34_17_n_4902, mul_34_17_n_4903, mul_34_17_n_4904, mul_34_17_n_4905,
     mul_34_17_n_4906, mul_34_17_n_4907, mul_34_17_n_4908, mul_34_17_n_4909,
     mul_34_17_n_4910, mul_34_17_n_4911, mul_34_17_n_4912, mul_34_17_n_4913,
     mul_34_17_n_4914, mul_34_17_n_4915, mul_34_17_n_4916, mul_34_17_n_4917,
     mul_34_17_n_4918, mul_34_17_n_4919, mul_34_17_n_4920, mul_34_17_n_4921,
     mul_34_17_n_4922, mul_34_17_n_4923, mul_34_17_n_4924, mul_34_17_n_4925,
     mul_34_17_n_4926, mul_34_17_n_4927, mul_34_17_n_4928, mul_34_17_n_4929,
     mul_34_17_n_4930, mul_34_17_n_4931, mul_34_17_n_4932, mul_34_17_n_4933,
     mul_34_17_n_4934, mul_34_17_n_4935, mul_34_17_n_4936, mul_34_17_n_4937,
     mul_34_17_n_4938, mul_34_17_n_4939, mul_34_17_n_4940, mul_34_17_n_4941,
     mul_34_17_n_4942, mul_34_17_n_4943, mul_34_17_n_4944, mul_34_17_n_4945,
     mul_34_17_n_4946, mul_34_17_n_4947, mul_34_17_n_4948, mul_34_17_n_4949,
     mul_34_17_n_4950, mul_34_17_n_4951, mul_34_17_n_4952, mul_34_17_n_4953,
     mul_34_17_n_4954, mul_34_17_n_4955, mul_34_17_n_4956, mul_34_17_n_4957,
     mul_34_17_n_4958, mul_34_17_n_4959, mul_34_17_n_4960, mul_34_17_n_4961,
     mul_34_17_n_4962, mul_34_17_n_4963, mul_34_17_n_4964, mul_34_17_n_4965,
     mul_34_17_n_4966, mul_34_17_n_4967, mul_34_17_n_4968, mul_34_17_n_4969,
     mul_34_17_n_4970, mul_34_17_n_4971, mul_34_17_n_4972, mul_34_17_n_4973,
     mul_34_17_n_4974, mul_34_17_n_4975, mul_34_17_n_4976, mul_34_17_n_4977,
     mul_34_17_n_4978, mul_34_17_n_4979, mul_34_17_n_4980, mul_34_17_n_4981,
     mul_34_17_n_4982, mul_34_17_n_4983, mul_34_17_n_4984, mul_34_17_n_4985,
     mul_34_17_n_4986, mul_34_17_n_4987, mul_34_17_n_4988, mul_34_17_n_4989,
     mul_34_17_n_4990, mul_34_17_n_4991, mul_34_17_n_4992, mul_34_17_n_4993,
     mul_34_17_n_4994, mul_34_17_n_4995, mul_34_17_n_4996, mul_34_17_n_4997,
     mul_34_17_n_4998, mul_34_17_n_4999, mul_34_17_n_5000, mul_34_17_n_5001,
     mul_34_17_n_5002, mul_34_17_n_5003, mul_34_17_n_5004, mul_34_17_n_5005,
     mul_34_17_n_5006, mul_34_17_n_5007, mul_34_17_n_5008, mul_34_17_n_5009,
     mul_34_17_n_5010, mul_34_17_n_5011, mul_34_17_n_5012, mul_34_17_n_5013,
     mul_34_17_n_5014, mul_34_17_n_5015, mul_34_17_n_5016, mul_34_17_n_5017,
     mul_34_17_n_5018, mul_34_17_n_5019, mul_34_17_n_5020, mul_34_17_n_5021,
     mul_34_17_n_5022, mul_34_17_n_5023, mul_34_17_n_5024, mul_34_17_n_5025,
     mul_34_17_n_5026, mul_34_17_n_5027, mul_34_17_n_5028, mul_34_17_n_5029,
     mul_34_17_n_5030, mul_34_17_n_5031, mul_34_17_n_5032, mul_34_17_n_5033,
     mul_34_17_n_5034, mul_34_17_n_5035, mul_34_17_n_5036, mul_34_17_n_5037,
     mul_34_17_n_5038, mul_34_17_n_5039, mul_34_17_n_5040, mul_34_17_n_5041,
     mul_34_17_n_5042, mul_34_17_n_5043, mul_34_17_n_5044, mul_34_17_n_5045,
     mul_34_17_n_5046, mul_34_17_n_5047, mul_34_17_n_5048, mul_34_17_n_5049,
     mul_34_17_n_5050, mul_34_17_n_5051, mul_34_17_n_5052, mul_34_17_n_5053,
     mul_34_17_n_5054, mul_34_17_n_5055, mul_34_17_n_5056, mul_34_17_n_5057,
     mul_34_17_n_5058, mul_34_17_n_5059, mul_34_17_n_5060, mul_34_17_n_5061,
     mul_34_17_n_5062, mul_34_17_n_5063, mul_34_17_n_5064, mul_34_17_n_5065,
     mul_34_17_n_5066, mul_34_17_n_5067, mul_34_17_n_5068, mul_34_17_n_5069,
     mul_34_17_n_5070, mul_34_17_n_5071, mul_34_17_n_5072, mul_34_17_n_5073,
     mul_34_17_n_5074, mul_34_17_n_5075, mul_34_17_n_5076, mul_34_17_n_5077,
     mul_34_17_n_5078, mul_34_17_n_5079, mul_34_17_n_5080, mul_34_17_n_5081,
     mul_34_17_n_5082, mul_34_17_n_5083, mul_34_17_n_5084, mul_34_17_n_5085,
     mul_34_17_n_5086, mul_34_17_n_5087, mul_34_17_n_5088, mul_34_17_n_5089,
     mul_34_17_n_5090, mul_34_17_n_5091, mul_34_17_n_5092, mul_34_17_n_5093,
     mul_34_17_n_5094, mul_34_17_n_5095, mul_34_17_n_5096, mul_34_17_n_5097,
     mul_34_17_n_5098, mul_34_17_n_5099, mul_34_17_n_5100, mul_34_17_n_5101,
     mul_34_17_n_5107, mul_34_17_n_5108, mul_34_17_n_5109, mul_34_17_n_5110,
     mul_34_17_n_5111, mul_34_17_n_5112, mul_34_17_n_5113, mul_34_17_n_5114,
     mul_34_17_n_5115, mul_34_17_n_5116, mul_34_17_n_5117, mul_34_17_n_5118,
     mul_34_17_n_5119, mul_34_17_n_5120, mul_34_17_n_5121, mul_34_17_n_5122,
     mul_34_17_n_5124, mul_34_17_n_5125, mul_34_17_n_5126, mul_34_17_n_5127,
     mul_34_17_n_5128, mul_34_17_n_5129, mul_34_17_n_5130, mul_34_17_n_5131,
     mul_34_17_n_5133, mul_34_17_n_5134, mul_34_17_n_5135, mul_34_17_n_5136,
     mul_34_17_n_5137, mul_34_17_n_5138, mul_34_17_n_5139, mul_34_17_n_5140,
     mul_34_17_n_5141, mul_34_17_n_5143, mul_34_17_n_5144, mul_34_17_n_5145,
     mul_34_17_n_5146, mul_34_17_n_5147, mul_34_17_n_5148, mul_34_17_n_5149,
     mul_34_17_n_5150, mul_34_17_n_5151, mul_34_17_n_5152, mul_34_17_n_5153,
     mul_34_17_n_5154, mul_34_17_n_5155, mul_34_17_n_5156, mul_34_17_n_5157,
     mul_34_17_n_5158, mul_34_17_n_5159, mul_34_17_n_5160, mul_34_17_n_5161,
     mul_34_17_n_5162, mul_34_17_n_5163, mul_34_17_n_5164, mul_34_17_n_5165,
     mul_34_17_n_5166, mul_34_17_n_5167, mul_34_17_n_5168, mul_34_17_n_5169,
     mul_34_17_n_5170, mul_34_17_n_5171, mul_34_17_n_5172, mul_34_17_n_5173,
     mul_34_17_n_5174, mul_34_17_n_5175, mul_34_17_n_5176, mul_34_17_n_5177,
     mul_34_17_n_5178, mul_34_17_n_5179, mul_34_17_n_5180, mul_34_17_n_5181,
     mul_34_17_n_5182, mul_34_17_n_5183, mul_34_17_n_5184, mul_34_17_n_5185,
     mul_34_17_n_5186, mul_34_17_n_5187, mul_34_17_n_5188, mul_34_17_n_5189,
     mul_34_17_n_5190, mul_34_17_n_5191, mul_34_17_n_5192, mul_34_17_n_5193,
     mul_34_17_n_5194, mul_34_17_n_5195, mul_34_17_n_5196, mul_34_17_n_5197,
     mul_34_17_n_5198, mul_34_17_n_5199, mul_34_17_n_5200, mul_34_17_n_5201,
     mul_34_17_n_5202, mul_34_17_n_5203, mul_34_17_n_5204, mul_34_17_n_5205,
     mul_34_17_n_5206, mul_34_17_n_5207, mul_34_17_n_5208, mul_34_17_n_5209,
     mul_34_17_n_5210, mul_34_17_n_5211, mul_34_17_n_5212, mul_34_17_n_5213,
     mul_34_17_n_5214, mul_34_17_n_5215, mul_34_17_n_5216, mul_34_17_n_5217,
     mul_34_17_n_5218, mul_34_17_n_5219, mul_34_17_n_5220, mul_34_17_n_5221,
     mul_34_17_n_5222, mul_34_17_n_5223, mul_34_17_n_5224, mul_34_17_n_5225,
     mul_34_17_n_5226, mul_34_17_n_5227, mul_34_17_n_5228, mul_34_17_n_5229,
     mul_34_17_n_5230, mul_34_17_n_5231, mul_34_17_n_5232, mul_34_17_n_5233,
     mul_34_17_n_5234, mul_34_17_n_5235, mul_34_17_n_5236, mul_34_17_n_5237,
     mul_34_17_n_5238, mul_34_17_n_5239, mul_34_17_n_5240, mul_34_17_n_5241,
     mul_34_17_n_5242, mul_34_17_n_5243, mul_34_17_n_5244, mul_34_17_n_5245,
     mul_34_17_n_5246, mul_34_17_n_5247, mul_34_17_n_5248, mul_34_17_n_5249,
     mul_34_17_n_5250, mul_34_17_n_5251, mul_34_17_n_5252, mul_34_17_n_5253,
     mul_34_17_n_5254, mul_34_17_n_5255, mul_34_17_n_5256, mul_34_17_n_5257,
     mul_34_17_n_5258, mul_34_17_n_5259, mul_34_17_n_5260, mul_34_17_n_5261,
     mul_34_17_n_5262, mul_34_17_n_5263, mul_34_17_n_5264, mul_34_17_n_5265,
     mul_34_17_n_5266, mul_34_17_n_5267, mul_34_17_n_5268, mul_34_17_n_5269,
     mul_34_17_n_5270, mul_34_17_n_5271, mul_34_17_n_5272, mul_34_17_n_5273,
     mul_34_17_n_5274, mul_34_17_n_5275, mul_34_17_n_5276, mul_34_17_n_5277,
     mul_34_17_n_5278, mul_34_17_n_5279, mul_34_17_n_5280, mul_34_17_n_5281,
     mul_34_17_n_5282, mul_34_17_n_5283, mul_34_17_n_5284, mul_34_17_n_5285,
     mul_34_17_n_5286, mul_34_17_n_5287, mul_34_17_n_5288, mul_34_17_n_5289,
     mul_34_17_n_5290, mul_34_17_n_5291, mul_34_17_n_5292, mul_34_17_n_5293,
     mul_34_17_n_5294, mul_34_17_n_5295, mul_34_17_n_5296, mul_34_17_n_5297,
     mul_34_17_n_5298, mul_34_17_n_5299, mul_34_17_n_5300, mul_34_17_n_5301,
     mul_34_17_n_5302, mul_34_17_n_5303, mul_34_17_n_5304, mul_34_17_n_5305,
     mul_34_17_n_5306, mul_34_17_n_5307, mul_34_17_n_5308, mul_34_17_n_5309,
     mul_34_17_n_5310, mul_34_17_n_5311, mul_34_17_n_5312, mul_34_17_n_5313,
     mul_34_17_n_5314, mul_34_17_n_5315, mul_34_17_n_5316, mul_34_17_n_5317,
     mul_34_17_n_5318, mul_34_17_n_5319, mul_34_17_n_5320, mul_34_17_n_5321,
     mul_34_17_n_5322, mul_34_17_n_5323, mul_34_17_n_5324, mul_34_17_n_5325,
     mul_34_17_n_5326, mul_34_17_n_5327, mul_34_17_n_5328, mul_34_17_n_5330,
     mul_34_17_n_5331, mul_34_17_n_5332, mul_34_17_n_5334, mul_34_17_n_5335,
     mul_34_17_n_5336, mul_34_17_n_5337, mul_34_17_n_5339, mul_34_17_n_5341,
     mul_34_17_n_5342, mul_34_17_n_5343, mul_34_17_n_5344, mul_34_17_n_5345,
     mul_34_17_n_5346, mul_34_17_n_5347, mul_34_17_n_5348, mul_34_17_n_5349,
     mul_34_17_n_5350, mul_34_17_n_5351, mul_34_17_n_5352, mul_34_17_n_5353,
     mul_34_17_n_5354, mul_34_17_n_5355, mul_34_17_n_5356, mul_34_17_n_5357,
     mul_34_17_n_5358, mul_34_17_n_5359, mul_34_17_n_5360, mul_34_17_n_5361,
     mul_34_17_n_5362, mul_34_17_n_5363, mul_34_17_n_5364, mul_34_17_n_5365,
     mul_34_17_n_5366, mul_34_17_n_5367, mul_34_17_n_5368, mul_34_17_n_5369,
     mul_34_17_n_5370, mul_34_17_n_5371, mul_34_17_n_5372, mul_34_17_n_5373,
     mul_34_17_n_5374, mul_34_17_n_5375, mul_34_17_n_5376, mul_34_17_n_5377,
     mul_34_17_n_5378, mul_34_17_n_5379, mul_34_17_n_5380, mul_34_17_n_5381,
     mul_34_17_n_5382, mul_34_17_n_5383, mul_34_17_n_5384, mul_34_17_n_5385,
     mul_34_17_n_5386, mul_34_17_n_5387, mul_34_17_n_5388, mul_34_17_n_5389,
     mul_34_17_n_5390, mul_34_17_n_5391, mul_34_17_n_5392, mul_34_17_n_5393,
     mul_34_17_n_5394, mul_34_17_n_5395, mul_34_17_n_5396, mul_34_17_n_5403,
     mul_34_17_n_5407, mul_34_17_n_5408, mul_34_17_n_5409, mul_34_17_n_5410,
     mul_34_17_n_5411, mul_34_17_n_5412, mul_34_17_n_5413, mul_34_17_n_5414,
     mul_34_17_n_5415, mul_34_17_n_5416, mul_34_17_n_5417, mul_34_17_n_5418,
     mul_34_17_n_5419, mul_34_17_n_5420, mul_34_17_n_5421, mul_34_17_n_5422,
     mul_34_17_n_5423, mul_34_17_n_5424, mul_34_17_n_5425, mul_34_17_n_5426,
     mul_34_17_n_5427, mul_34_17_n_5428, mul_34_17_n_5429, mul_34_17_n_5430,
     mul_34_17_n_5431, mul_34_17_n_5432, mul_34_17_n_5433, mul_34_17_n_5434,
     mul_34_17_n_5435, mul_34_17_n_5436, mul_34_17_n_5437, mul_34_17_n_5438,
     mul_34_17_n_5439, mul_34_17_n_5440, mul_34_17_n_5441, mul_34_17_n_5442,
     mul_34_17_n_5443, mul_34_17_n_5444, mul_34_17_n_5445, mul_34_17_n_5446,
     mul_34_17_n_5447, mul_34_17_n_5448, mul_34_17_n_5449, mul_34_17_n_5450,
     mul_34_17_n_5451, mul_34_17_n_5452, mul_34_17_n_5453, mul_34_17_n_5454,
     mul_34_17_n_5455, mul_34_17_n_5456, mul_34_17_n_5457, mul_34_17_n_5458,
     mul_34_17_n_5459, mul_34_17_n_5460, mul_34_17_n_5461, mul_34_17_n_5462,
     mul_34_17_n_5463, mul_34_17_n_5464, mul_34_17_n_5465, mul_34_17_n_5466,
     mul_34_17_n_5467, mul_34_17_n_5468, mul_34_17_n_5469, mul_34_17_n_5470,
     mul_34_17_n_5471, mul_34_17_n_5472, mul_34_17_n_5473, mul_34_17_n_5474,
     mul_34_17_n_5475, mul_34_17_n_5476, mul_34_17_n_5477, mul_34_17_n_5478,
     mul_34_17_n_5479, mul_34_17_n_5480, mul_34_17_n_5481, mul_34_17_n_5482,
     mul_34_17_n_5483, mul_34_17_n_5484, mul_34_17_n_5485, mul_34_17_n_5486,
     mul_34_17_n_5487, mul_34_17_n_5488, mul_34_17_n_5489, mul_34_17_n_5490,
     mul_34_17_n_5491, mul_34_17_n_5492, mul_34_17_n_5493, mul_34_17_n_5494,
     mul_34_17_n_5495, mul_34_17_n_5496, mul_34_17_n_5497, mul_34_17_n_5498,
     mul_34_17_n_5499, mul_34_17_n_5500, mul_34_17_n_5501, mul_34_17_n_5502,
     mul_34_17_n_5503, mul_34_17_n_5504, mul_34_17_n_5505, mul_34_17_n_5506,
     mul_34_17_n_5507, mul_34_17_n_5508, mul_34_17_n_5509, mul_34_17_n_5510,
     mul_34_17_n_5511, mul_34_17_n_5512, mul_34_17_n_5513, mul_34_17_n_5514,
     mul_34_17_n_5515, mul_34_17_n_5516, mul_34_17_n_5517, mul_34_17_n_5518,
     mul_34_17_n_5519, mul_34_17_n_5520, mul_34_17_n_5521, mul_34_17_n_5522,
     mul_34_17_n_5523, mul_34_17_n_5524, mul_34_17_n_5525, mul_34_17_n_5526,
     mul_34_17_n_5527, mul_34_17_n_5528, mul_34_17_n_5529, mul_34_17_n_5530,
     mul_34_17_n_5531, mul_34_17_n_5532, mul_34_17_n_5533, mul_34_17_n_5534,
     mul_34_17_n_5535, mul_34_17_n_5536, mul_34_17_n_5537, mul_34_17_n_5538,
     mul_34_17_n_5539, mul_34_17_n_5540, mul_34_17_n_5541, mul_34_17_n_5542,
     mul_34_17_n_5543, mul_34_17_n_5544, mul_34_17_n_5545, mul_34_17_n_5546,
     mul_34_17_n_5547, mul_34_17_n_5548, mul_34_17_n_5549, mul_34_17_n_5550,
     mul_34_17_n_5551, mul_34_17_n_5552, mul_34_17_n_5553, mul_34_17_n_5554,
     mul_34_17_n_5555, mul_34_17_n_5556, mul_34_17_n_5557, mul_34_17_n_5558,
     mul_34_17_n_5559, mul_34_17_n_5560, mul_34_17_n_5561, mul_34_17_n_5562,
     mul_34_17_n_5563, mul_34_17_n_5564, mul_34_17_n_5565, mul_34_17_n_5566,
     mul_34_17_n_5567, mul_34_17_n_5568, mul_34_17_n_5569, mul_34_17_n_5570,
     mul_34_17_n_5571, mul_34_17_n_5572, mul_34_17_n_5573, mul_34_17_n_5574,
     mul_34_17_n_5575, mul_34_17_n_5576, mul_34_17_n_5577, mul_34_17_n_5578,
     mul_34_17_n_5579, mul_34_17_n_5580, mul_34_17_n_5581, mul_34_17_n_5582,
     mul_34_17_n_5583, mul_34_17_n_5584, mul_34_17_n_5585, mul_34_17_n_5586,
     mul_34_17_n_5587, mul_34_17_n_5588, mul_34_17_n_5589, mul_34_17_n_5590,
     mul_34_17_n_5591, mul_34_17_n_5592, mul_34_17_n_5593, mul_34_17_n_5594,
     mul_34_17_n_5595, mul_34_17_n_5596, mul_34_17_n_5597, mul_34_17_n_5598,
     mul_34_17_n_5599, mul_34_17_n_5600, mul_34_17_n_5601, mul_34_17_n_5602,
     mul_34_17_n_5603, mul_34_17_n_5604, mul_34_17_n_5605, mul_34_17_n_5606,
     mul_34_17_n_5607, mul_34_17_n_5608, mul_34_17_n_5609, mul_34_17_n_5610,
     mul_34_17_n_5611, mul_34_17_n_5612, mul_34_17_n_5613, mul_34_17_n_5614,
     mul_34_17_n_5615, mul_34_17_n_5616, mul_34_17_n_5617, mul_34_17_n_5618,
     mul_34_17_n_5619, mul_34_17_n_5620, mul_34_17_n_5621, mul_34_17_n_5622,
     mul_34_17_n_5623, mul_34_17_n_5624, mul_34_17_n_5625, mul_34_17_n_5626,
     mul_34_17_n_5627, mul_34_17_n_5628, mul_34_17_n_5629, mul_34_17_n_5630,
     mul_34_17_n_5631, mul_34_17_n_5632, mul_34_17_n_5633, mul_34_17_n_5634,
     mul_34_17_n_5635, mul_34_17_n_5636, mul_34_17_n_5637, mul_34_17_n_5638,
     mul_34_17_n_5639, mul_34_17_n_5640, mul_34_17_n_5641, mul_34_17_n_5642,
     mul_34_17_n_5643, mul_34_17_n_5644, mul_34_17_n_5645, mul_34_17_n_5646,
     mul_34_17_n_5647, mul_34_17_n_5648, mul_34_17_n_5649, mul_34_17_n_5650,
     mul_34_17_n_5651, mul_34_17_n_5652, mul_34_17_n_5653, mul_34_17_n_5654,
     mul_34_17_n_5655, mul_34_17_n_5656, mul_34_17_n_5657, mul_34_17_n_5658,
     mul_34_17_n_5659, mul_34_17_n_5660, mul_34_17_n_5661, mul_34_17_n_5662,
     mul_34_17_n_5663, mul_34_17_n_5664, mul_34_17_n_5665, mul_34_17_n_5666,
     mul_34_17_n_5667, mul_34_17_n_5668, mul_34_17_n_5669, mul_34_17_n_5670,
     mul_34_17_n_5671, mul_34_17_n_5672, mul_34_17_n_5673, mul_34_17_n_5674,
     mul_34_17_n_5675, mul_34_17_n_5676, mul_34_17_n_5677, mul_34_17_n_5678,
     mul_34_17_n_5679, mul_34_17_n_5680, mul_34_17_n_5681, mul_34_17_n_5682,
     mul_34_17_n_5683, mul_34_17_n_5684, mul_34_17_n_5685, mul_34_17_n_5686,
     mul_34_17_n_5687, mul_34_17_n_5688, mul_34_17_n_5689, mul_34_17_n_5690,
     mul_34_17_n_5691, mul_34_17_n_5692, mul_34_17_n_5693, mul_34_17_n_5694,
     mul_34_17_n_5695, mul_34_17_n_5696, mul_34_17_n_5697, mul_34_17_n_5698,
     mul_34_17_n_5699, mul_34_17_n_5700, mul_34_17_n_5701, mul_34_17_n_5702,
     mul_34_17_n_5703, mul_34_17_n_5704, mul_34_17_n_5705, mul_34_17_n_5706,
     mul_34_17_n_5707, mul_34_17_n_5708, mul_34_17_n_5709, mul_34_17_n_5710,
     mul_34_17_n_5711, mul_34_17_n_5712, mul_34_17_n_5713, mul_34_17_n_5714,
     mul_34_17_n_5715, mul_34_17_n_5716, mul_34_17_n_5717, mul_34_17_n_5718,
     mul_34_17_n_5719, mul_34_17_n_5720, mul_34_17_n_5721, mul_34_17_n_5722,
     mul_34_17_n_5723, mul_34_17_n_5724, mul_34_17_n_5725, mul_34_17_n_5726,
     mul_34_17_n_5727, mul_34_17_n_5728, mul_34_17_n_5729, mul_34_17_n_5730,
     mul_34_17_n_5731, mul_34_17_n_5732, mul_34_17_n_5733, mul_34_17_n_5734,
     mul_34_17_n_5735, mul_34_17_n_5736, mul_34_17_n_5737, mul_34_17_n_5738,
     mul_34_17_n_5739, mul_34_17_n_5740, mul_34_17_n_5741, mul_34_17_n_5742,
     mul_34_17_n_5743, mul_34_17_n_5744, mul_34_17_n_5745, mul_34_17_n_5746,
     mul_34_17_n_5747, mul_34_17_n_5748, mul_34_17_n_5749, mul_34_17_n_5750,
     mul_34_17_n_5751, mul_34_17_n_5752, mul_34_17_n_5753, mul_34_17_n_5754,
     mul_34_17_n_5755, mul_34_17_n_5756, mul_34_17_n_5757, mul_34_17_n_5758,
     mul_34_17_n_5759, mul_34_17_n_5760, mul_34_17_n_5761, mul_34_17_n_5762,
     mul_34_17_n_5763, mul_34_17_n_5764, mul_34_17_n_5765, mul_34_17_n_5766,
     mul_34_17_n_5767, mul_34_17_n_5768, mul_34_17_n_5769, mul_34_17_n_5770,
     mul_34_17_n_5771, mul_34_17_n_5772, mul_34_17_n_5773, mul_34_17_n_5774,
     mul_34_17_n_5775, mul_34_17_n_5776, mul_34_17_n_5777, mul_34_17_n_5778,
     mul_34_17_n_5779, mul_34_17_n_5780, mul_34_17_n_5781, mul_34_17_n_5782,
     mul_34_17_n_5783, mul_34_17_n_5784, mul_34_17_n_5785, mul_34_17_n_5786,
     mul_34_17_n_5787, mul_34_17_n_5788, mul_34_17_n_5789, mul_34_17_n_5790,
     mul_34_17_n_5791, mul_34_17_n_5792, mul_34_17_n_5793, mul_34_17_n_5794,
     mul_34_17_n_5795, mul_34_17_n_5796, mul_34_17_n_5797, mul_34_17_n_5798,
     mul_34_17_n_5799, mul_34_17_n_5800, mul_34_17_n_5801, mul_34_17_n_5802,
     mul_34_17_n_5803, mul_34_17_n_5804, mul_34_17_n_5805, mul_34_17_n_5806,
     mul_34_17_n_5807, mul_34_17_n_5808, mul_34_17_n_5809, mul_34_17_n_5810,
     mul_34_17_n_5811, mul_34_17_n_5812, mul_34_17_n_5813, mul_34_17_n_5814,
     mul_34_17_n_5816, mul_34_17_n_5817, mul_34_17_n_5818, mul_34_17_n_5819,
     mul_34_17_n_5820, mul_34_17_n_5821, mul_34_17_n_5822, mul_34_17_n_5823,
     mul_34_17_n_5824, mul_34_17_n_5825, mul_34_17_n_5826, mul_34_17_n_5827,
     mul_34_17_n_5828, mul_34_17_n_5829, mul_34_17_n_5830, mul_34_17_n_5831,
     mul_34_17_n_5832, mul_34_17_n_5833, mul_34_17_n_5834, mul_34_17_n_5835,
     mul_34_17_n_5836, mul_34_17_n_5838, mul_34_17_n_5839, mul_34_17_n_5840,
     mul_34_17_n_5841, mul_34_17_n_5842, mul_34_17_n_5843, mul_34_17_n_5844,
     mul_34_17_n_5845, mul_34_17_n_5846, mul_34_17_n_5847, mul_34_17_n_5848,
     mul_34_17_n_5849, mul_34_17_n_5850, mul_34_17_n_5851, mul_34_17_n_5852,
     mul_34_17_n_5853, mul_34_17_n_5854, mul_34_17_n_5855, mul_34_17_n_5856,
     mul_34_17_n_5857, mul_34_17_n_5858, mul_34_17_n_5859, mul_34_17_n_5860,
     mul_34_17_n_5861, mul_34_17_n_5862, mul_34_17_n_5863, mul_34_17_n_5864,
     mul_34_17_n_5865, mul_34_17_n_5866, mul_34_17_n_5867, mul_34_17_n_5868,
     mul_34_17_n_5869, mul_34_17_n_5870, mul_34_17_n_5871, mul_34_17_n_5872,
     mul_34_17_n_5874, mul_34_17_n_5875, mul_34_17_n_5876, mul_34_17_n_5877,
     mul_34_17_n_5878, mul_34_17_n_5879, mul_34_17_n_5880, mul_34_17_n_5881,
     mul_34_17_n_5882, mul_34_17_n_5883, mul_34_17_n_5884, mul_34_17_n_5885,
     mul_34_17_n_5886, mul_34_17_n_5887, mul_34_17_n_5888, mul_34_17_n_5889,
     mul_34_17_n_5890, mul_34_17_n_5891, mul_34_17_n_5892, mul_34_17_n_5893,
     mul_34_17_n_5894, mul_34_17_n_5895, mul_34_17_n_5896, mul_34_17_n_5897,
     mul_34_17_n_5898, mul_34_17_n_5899, mul_34_17_n_5900, mul_34_17_n_5901,
     mul_34_17_n_5902, mul_34_17_n_5903, mul_34_17_n_5904, mul_34_17_n_5905,
     mul_34_17_n_5906, mul_34_17_n_5907, mul_34_17_n_5908, mul_34_17_n_5909,
     mul_34_17_n_5910, mul_34_17_n_5911, mul_34_17_n_5912, mul_34_17_n_5913,
     mul_34_17_n_5914, mul_34_17_n_5915, mul_34_17_n_5916, mul_34_17_n_5917,
     mul_34_17_n_5918, mul_34_17_n_5919, mul_34_17_n_5920, mul_34_17_n_5921,
     mul_34_17_n_5922, mul_34_17_n_5923, mul_34_17_n_5924, mul_34_17_n_5925,
     mul_34_17_n_5926, mul_34_17_n_5927, mul_34_17_n_5928, mul_34_17_n_5929,
     mul_34_17_n_5930, mul_34_17_n_5931, mul_34_17_n_5932, mul_34_17_n_5933,
     mul_34_17_n_5934, mul_34_17_n_5935, mul_34_17_n_5936, mul_34_17_n_5937,
     mul_34_17_n_5938, mul_34_17_n_5939, mul_34_17_n_5940, mul_34_17_n_5941,
     mul_34_17_n_5942, mul_34_17_n_5943, mul_34_17_n_5944, mul_34_17_n_5945,
     mul_34_17_n_5946, mul_34_17_n_5947, mul_34_17_n_5948, mul_34_17_n_5949,
     mul_34_17_n_5950, mul_34_17_n_5951, mul_34_17_n_5952, mul_34_17_n_5953,
     mul_34_17_n_5954, mul_34_17_n_5955, mul_34_17_n_5956, mul_34_17_n_5957,
     mul_34_17_n_5958, mul_34_17_n_5959, mul_34_17_n_5960, mul_34_17_n_5961,
     mul_34_17_n_5962, mul_34_17_n_5963, mul_34_17_n_5964, mul_34_17_n_5965,
     mul_34_17_n_5966, mul_34_17_n_5967, mul_34_17_n_5968, mul_34_17_n_5969,
     mul_34_17_n_5970, mul_34_17_n_5971, mul_34_17_n_5972, mul_34_17_n_5973,
     mul_34_17_n_5974, mul_34_17_n_5975, mul_34_17_n_5976, mul_34_17_n_5977,
     mul_34_17_n_5978, mul_34_17_n_5979, mul_34_17_n_5980, mul_34_17_n_5981,
     mul_34_17_n_5982, mul_34_17_n_5983, mul_34_17_n_5984, mul_34_17_n_5985,
     mul_34_17_n_5986, mul_34_17_n_5987, mul_34_17_n_5988, mul_34_17_n_5989,
     mul_34_17_n_5990, mul_34_17_n_5991, mul_34_17_n_5992, mul_34_17_n_5993,
     mul_34_17_n_5994, mul_34_17_n_5995, mul_34_17_n_5996, mul_34_17_n_5997,
     mul_34_17_n_5998, mul_34_17_n_5999, mul_34_17_n_6000, mul_34_17_n_6001,
     mul_34_17_n_6002, mul_34_17_n_6003, mul_34_17_n_6004, mul_34_17_n_6005,
     mul_34_17_n_6006, mul_34_17_n_6007, mul_34_17_n_6008, mul_34_17_n_6009,
     mul_34_17_n_6010, mul_34_17_n_6011, mul_34_17_n_6012, mul_34_17_n_6013,
     mul_34_17_n_6014, mul_34_17_n_6015, mul_34_17_n_6016, mul_34_17_n_6017,
     mul_34_17_n_6018, mul_34_17_n_6019, mul_34_17_n_6020, mul_34_17_n_6021,
     mul_34_17_n_6022, mul_34_17_n_6023, mul_34_17_n_6024, mul_34_17_n_6025,
     mul_34_17_n_6026, mul_34_17_n_6027, mul_34_17_n_6028, mul_34_17_n_6029,
     mul_34_17_n_6030, mul_34_17_n_6031, mul_34_17_n_6032, mul_34_17_n_6033,
     mul_34_17_n_6034, mul_34_17_n_6035, mul_34_17_n_6036, mul_34_17_n_6037,
     mul_34_17_n_6038, mul_34_17_n_6039, mul_34_17_n_6040, mul_34_17_n_6041,
     mul_34_17_n_6042, mul_34_17_n_6043, mul_34_17_n_6044, mul_34_17_n_6045,
     mul_34_17_n_6046, mul_34_17_n_6047, mul_34_17_n_6048, mul_34_17_n_6049,
     mul_34_17_n_6050, mul_34_17_n_6051, mul_34_17_n_6052, mul_34_17_n_6053,
     mul_34_17_n_6054, mul_34_17_n_6055, mul_34_17_n_6056, mul_34_17_n_6057,
     mul_34_17_n_6058, mul_34_17_n_6059, mul_34_17_n_6060, mul_34_17_n_6061,
     mul_34_17_n_6062, mul_34_17_n_6063, mul_34_17_n_6064, mul_34_17_n_6065,
     mul_34_17_n_6066, mul_34_17_n_6067, mul_34_17_n_6068, mul_34_17_n_6069,
     mul_34_17_n_6070, mul_34_17_n_6071, mul_34_17_n_6072, mul_34_17_n_6073,
     mul_34_17_n_6074, mul_34_17_n_6075, mul_34_17_n_6076, mul_34_17_n_6077,
     mul_34_17_n_6078, mul_34_17_n_6079, mul_34_17_n_6080, mul_34_17_n_6081,
     mul_34_17_n_6082, mul_34_17_n_6083, mul_34_17_n_6084, mul_34_17_n_6085,
     mul_34_17_n_6086, mul_34_17_n_6087, mul_34_17_n_6088, mul_34_17_n_6089,
     mul_34_17_n_6090, mul_34_17_n_6091, mul_34_17_n_6092, mul_34_17_n_6093,
     mul_34_17_n_6094, mul_34_17_n_6095, mul_34_17_n_6096, mul_34_17_n_6097,
     mul_34_17_n_6098, mul_34_17_n_6099, mul_34_17_n_6100, mul_34_17_n_6101,
     mul_34_17_n_6102, mul_34_17_n_6103, mul_34_17_n_6104, mul_34_17_n_6105,
     mul_34_17_n_6106, mul_34_17_n_6107, mul_34_17_n_6108, mul_34_17_n_6109,
     mul_34_17_n_6110, mul_34_17_n_6111, mul_34_17_n_6112, mul_34_17_n_6113,
     mul_34_17_n_6114, mul_34_17_n_6115, mul_34_17_n_6116, mul_34_17_n_6117,
     mul_34_17_n_6118, mul_34_17_n_6119, mul_34_17_n_6120, mul_34_17_n_6121,
     mul_34_17_n_6122, mul_34_17_n_6123, mul_34_17_n_6124, mul_34_17_n_6125,
     mul_34_17_n_6126, mul_34_17_n_6127, mul_34_17_n_6128, mul_34_17_n_6129,
     mul_34_17_n_6130, mul_34_17_n_6131, mul_34_17_n_6132, mul_34_17_n_6133,
     mul_34_17_n_6134, mul_34_17_n_6135, mul_34_17_n_6136, mul_34_17_n_6137,
     mul_34_17_n_6138, mul_34_17_n_6139, mul_34_17_n_6140, mul_34_17_n_6141,
     mul_34_17_n_6142, mul_34_17_n_6143, mul_34_17_n_6144, mul_34_17_n_6145,
     mul_34_17_n_6146, mul_34_17_n_6147, mul_34_17_n_6152, mul_34_17_n_6153,
     mul_34_17_n_6154, mul_34_17_n_6155, mul_34_17_n_6156, mul_34_17_n_6158,
     mul_34_17_n_6159, mul_34_17_n_6160, mul_34_17_n_6161, mul_34_17_n_6162,
     mul_34_17_n_6163, mul_34_17_n_6164, mul_34_17_n_6165, mul_34_17_n_6166,
     mul_34_17_n_6167, mul_34_17_n_6168, mul_34_17_n_6169, mul_34_17_n_6170,
     mul_34_17_n_6171, mul_34_17_n_6172, mul_34_17_n_6173, mul_34_17_n_6174,
     mul_34_17_n_6175, mul_34_17_n_6176, mul_34_17_n_6177, mul_34_17_n_6178,
     mul_34_17_n_6179, mul_34_17_n_6181, mul_34_17_n_6182, mul_34_17_n_6183,
     mul_34_17_n_6184, mul_34_17_n_6185, mul_34_17_n_6186, mul_34_17_n_6188,
     mul_34_17_n_6189, mul_34_17_n_6190, mul_34_17_n_6191, mul_34_17_n_6192,
     mul_34_17_n_6193, mul_34_17_n_6194, mul_34_17_n_6195, mul_34_17_n_6196,
     mul_34_17_n_6197, mul_34_17_n_6198, mul_34_17_n_6199, mul_34_17_n_6200,
     mul_34_17_n_6201, mul_34_17_n_6202, mul_34_17_n_6203, mul_34_17_n_6204,
     mul_34_17_n_6205, mul_34_17_n_6206, mul_34_17_n_6208, mul_34_17_n_6209,
     mul_34_17_n_6210, mul_34_17_n_6211, mul_34_17_n_6212, mul_34_17_n_6213,
     mul_34_17_n_6214, mul_34_17_n_6215, mul_34_17_n_6216, mul_34_17_n_6217,
     mul_34_17_n_6218, mul_34_17_n_6219, mul_34_17_n_6220, mul_34_17_n_6221,
     mul_34_17_n_6222, mul_34_17_n_6223, mul_34_17_n_6224, mul_34_17_n_6225,
     mul_34_17_n_6226, mul_34_17_n_6227, mul_34_17_n_6228, mul_34_17_n_6229,
     mul_34_17_n_6230, mul_34_17_n_6231, mul_34_17_n_6232, mul_34_17_n_6233,
     mul_34_17_n_6234, mul_34_17_n_6235, mul_34_17_n_6236, mul_34_17_n_6237,
     mul_34_17_n_6239, mul_34_17_n_6240, mul_34_17_n_6241, mul_34_17_n_6242,
     mul_34_17_n_6243, mul_34_17_n_6244, mul_34_17_n_6245, mul_34_17_n_6246,
     mul_34_17_n_6247, mul_34_17_n_6248, mul_34_17_n_6249, mul_34_17_n_6250,
     mul_34_17_n_6251, mul_34_17_n_6252, mul_34_17_n_6253, mul_34_17_n_6254,
     mul_34_17_n_6255, mul_34_17_n_6256, mul_34_17_n_6259, mul_34_17_n_6260,
     mul_34_17_n_6261, mul_34_17_n_6262, mul_34_17_n_6265, mul_34_17_n_6266,
     mul_34_17_n_6267, mul_34_17_n_6268, mul_34_17_n_6269, mul_34_17_n_6270,
     mul_34_17_n_6271, mul_34_17_n_6273, mul_34_17_n_6275, mul_34_17_n_6277,
     mul_34_17_n_6278, mul_34_17_n_6280, mul_34_17_n_6281, mul_34_17_n_6282,
     mul_34_17_n_6283, mul_34_17_n_6284, mul_34_17_n_6285, mul_34_17_n_6286,
     mul_34_17_n_6287, mul_34_17_n_6289, mul_34_17_n_6290, mul_34_17_n_6291,
     mul_34_17_n_6294, mul_34_17_n_6295, mul_34_17_n_6296, mul_34_17_n_6297,
     mul_34_17_n_6298, mul_34_17_n_6299, mul_34_17_n_6300, mul_34_17_n_6301,
     mul_34_17_n_6302, mul_34_17_n_6303, mul_34_17_n_6304, mul_34_17_n_6305,
     mul_34_17_n_6306, mul_34_17_n_6307, mul_34_17_n_6308, mul_34_17_n_6309,
     mul_34_17_n_6311, mul_34_17_n_6312, mul_34_17_n_6313, mul_34_17_n_6315,
     mul_34_17_n_6316, mul_34_17_n_6317, mul_34_17_n_6318, mul_34_17_n_6319,
     mul_34_17_n_6320, mul_34_17_n_6322, mul_34_17_n_6323, mul_34_17_n_6324,
     mul_34_17_n_6325, mul_34_17_n_6326, mul_34_17_n_6327, mul_34_17_n_6328,
     mul_34_17_n_6329, mul_34_17_n_6330, mul_34_17_n_6331, mul_34_17_n_6332,
     mul_34_17_n_6333, mul_34_17_n_6334, mul_34_17_n_6335, mul_34_17_n_6336,
     mul_34_17_n_6338, mul_34_17_n_6340, mul_34_17_n_6341, mul_34_17_n_6342,
     mul_34_17_n_6343, mul_34_17_n_6344, mul_34_17_n_6345, mul_34_17_n_6346,
     mul_34_17_n_6347, mul_34_17_n_6348, mul_34_17_n_6349, mul_34_17_n_6350,
     mul_34_17_n_6351, mul_34_17_n_6352, mul_34_17_n_6353, mul_34_17_n_6354,
     mul_34_17_n_6355, mul_34_17_n_6356, mul_34_17_n_6357, mul_34_17_n_6358,
     mul_34_17_n_6360, mul_34_17_n_6361, mul_34_17_n_6362, mul_34_17_n_6363,
     mul_34_17_n_6364, mul_34_17_n_6365, mul_34_17_n_6366, mul_34_17_n_6367,
     mul_34_17_n_6368, mul_34_17_n_6369, mul_34_17_n_6370, mul_34_17_n_6371,
     mul_34_17_n_6373, mul_34_17_n_6374, mul_34_17_n_6375, mul_34_17_n_6376,
     mul_34_17_n_6377, mul_34_17_n_6379, mul_34_17_n_6380, mul_34_17_n_6381,
     mul_34_17_n_6382, mul_34_17_n_6384, mul_34_17_n_6385, mul_34_17_n_6387,
     mul_34_17_n_6388, mul_34_17_n_6389, mul_34_17_n_6390, mul_34_17_n_6391,
     mul_34_17_n_6392, mul_34_17_n_6393, mul_34_17_n_6394, mul_34_17_n_6395,
     mul_34_17_n_6396, mul_34_17_n_6397, mul_34_17_n_6398, mul_34_17_n_6399,
     mul_34_17_n_6400, mul_34_17_n_6401, mul_34_17_n_6402, mul_34_17_n_6403,
     mul_34_17_n_6404, mul_34_17_n_6405, mul_34_17_n_6406, mul_34_17_n_6407,
     mul_34_17_n_6408, mul_34_17_n_6409, mul_34_17_n_6411, mul_34_17_n_6412,
     mul_34_17_n_6413, mul_34_17_n_6414, mul_34_17_n_6415, mul_34_17_n_6416,
     mul_34_17_n_6417, mul_34_17_n_6418, mul_34_17_n_6419, mul_34_17_n_6420,
     mul_34_17_n_6421, mul_34_17_n_6422, mul_34_17_n_6423, mul_34_17_n_6424,
     mul_34_17_n_6425, mul_34_17_n_6426, mul_34_17_n_6427, mul_34_17_n_6428,
     mul_34_17_n_6429, mul_34_17_n_6430, mul_34_17_n_6431, mul_34_17_n_6432,
     mul_34_17_n_6433, mul_34_17_n_6434, mul_34_17_n_6435, mul_34_17_n_6436,
     mul_34_17_n_6437, mul_34_17_n_6438, mul_34_17_n_6439, mul_34_17_n_6440,
     mul_34_17_n_6441, mul_34_17_n_6442, mul_34_17_n_6443, mul_34_17_n_6444,
     mul_34_17_n_6445, mul_34_17_n_6446, mul_34_17_n_6447, mul_34_17_n_6448,
     mul_34_17_n_6449, mul_34_17_n_6450, mul_34_17_n_6451, mul_34_17_n_6452,
     mul_34_17_n_6454, mul_34_17_n_6455, mul_34_17_n_6456, mul_34_17_n_6457,
     mul_34_17_n_6458, mul_34_17_n_6459, mul_34_17_n_6460, mul_34_17_n_6461,
     mul_34_17_n_6462, mul_34_17_n_6464, mul_34_17_n_6465, mul_34_17_n_6466,
     mul_34_17_n_6467, mul_34_17_n_6469, mul_34_17_n_6471, mul_34_17_n_6472,
     mul_34_17_n_6474, mul_34_17_n_6476, mul_34_17_n_6477, mul_34_17_n_6478,
     mul_34_17_n_6479, mul_34_17_n_6480, mul_34_17_n_6481, mul_34_17_n_6482,
     mul_34_17_n_6483, mul_34_17_n_6484, mul_34_17_n_6486, mul_34_17_n_6487,
     mul_34_17_n_6488, mul_34_17_n_6489, mul_34_17_n_6490, mul_34_17_n_6491,
     mul_34_17_n_6492, mul_34_17_n_6493, mul_34_17_n_6495, mul_34_17_n_6497,
     mul_34_17_n_6498, mul_34_17_n_6499, mul_34_17_n_6500, mul_34_17_n_6501,
     mul_34_17_n_6502, mul_34_17_n_6503, mul_34_17_n_6504, mul_34_17_n_6505,
     mul_34_17_n_6506, mul_34_17_n_6507, mul_34_17_n_6508, mul_34_17_n_6509,
     mul_34_17_n_6510, mul_34_17_n_6511, mul_34_17_n_6512, mul_34_17_n_6513,
     mul_34_17_n_6514, mul_34_17_n_6516, mul_34_17_n_6517, mul_34_17_n_6518,
     mul_34_17_n_6519, mul_34_17_n_6520, mul_34_17_n_6521, mul_34_17_n_6522,
     mul_34_17_n_6523, mul_34_17_n_6524, mul_34_17_n_6525, mul_34_17_n_6526,
     mul_34_17_n_6527, mul_34_17_n_6528, mul_34_17_n_6529, mul_34_17_n_6530,
     mul_34_17_n_6531, mul_34_17_n_6532, mul_34_17_n_6533, mul_34_17_n_6534,
     mul_34_17_n_6535, mul_34_17_n_6536, mul_34_17_n_6537, mul_34_17_n_6538,
     mul_34_17_n_6539, mul_34_17_n_6540, mul_34_17_n_6541, mul_34_17_n_6542,
     mul_34_17_n_6543, mul_34_17_n_6544, mul_34_17_n_6545, mul_34_17_n_6546,
     mul_34_17_n_6547, mul_34_17_n_6548, mul_34_17_n_6550, mul_34_17_n_6552,
     mul_34_17_n_6553, mul_34_17_n_6554, mul_34_17_n_6556, mul_34_17_n_6557,
     mul_34_17_n_6559, mul_34_17_n_6560, mul_34_17_n_6561, mul_34_17_n_6562,
     mul_34_17_n_6563, mul_34_17_n_6564, mul_34_17_n_6565, mul_34_17_n_6566,
     mul_34_17_n_6567, mul_34_17_n_6568, mul_34_17_n_6570, mul_34_17_n_6571,
     mul_34_17_n_6572, mul_34_17_n_6573, mul_34_17_n_6574, mul_34_17_n_6575,
     mul_34_17_n_6576, mul_34_17_n_6577, mul_34_17_n_6579, mul_34_17_n_6581,
     mul_34_17_n_6584, mul_34_17_n_6585, mul_34_17_n_6586, mul_34_17_n_6588,
     mul_34_17_n_6589, mul_34_17_n_6590, mul_34_17_n_6591, mul_34_17_n_6593,
     mul_34_17_n_6594, mul_34_17_n_6595, mul_34_17_n_6596, mul_34_17_n_6597,
     mul_34_17_n_6598, mul_34_17_n_6599, mul_34_17_n_6600, mul_34_17_n_6601,
     mul_34_17_n_6602, mul_34_17_n_6603, mul_34_17_n_6604, mul_34_17_n_6605,
     mul_34_17_n_6606, mul_34_17_n_6607, mul_34_17_n_6608, mul_34_17_n_6609,
     mul_34_17_n_6610, mul_34_17_n_6611, mul_34_17_n_6613, mul_34_17_n_6614,
     mul_34_17_n_6615, mul_34_17_n_6616, mul_34_17_n_6617, mul_34_17_n_6618,
     mul_34_17_n_6619, mul_34_17_n_6620, mul_34_17_n_6621, mul_34_17_n_6622,
     mul_34_17_n_6623, mul_34_17_n_6624, mul_34_17_n_6625, mul_34_17_n_6626,
     mul_34_17_n_6627, mul_34_17_n_6628, mul_34_17_n_6629, mul_34_17_n_6630,
     mul_34_17_n_6631, mul_34_17_n_6632, mul_34_17_n_6633, mul_34_17_n_6634,
     mul_34_17_n_6635, mul_34_17_n_6636, mul_34_17_n_6637, mul_34_17_n_6638,
     mul_34_17_n_6639, mul_34_17_n_6640, mul_34_17_n_6641, mul_34_17_n_6642,
     mul_34_17_n_6643, mul_34_17_n_6644, mul_34_17_n_6645, mul_34_17_n_6646,
     mul_34_17_n_6647, mul_34_17_n_6648, mul_34_17_n_6649, mul_34_17_n_6650,
     mul_34_17_n_6652, mul_34_17_n_6653, mul_34_17_n_6654, mul_34_17_n_6655,
     mul_34_17_n_6657, mul_34_17_n_6659, mul_34_17_n_6660, mul_34_17_n_6661,
     mul_34_17_n_6662, mul_34_17_n_6663, mul_34_17_n_6664, mul_34_17_n_6665,
     mul_34_17_n_6666, mul_34_17_n_6667, mul_34_17_n_6668, mul_34_17_n_6670,
     mul_34_17_n_6671, mul_34_17_n_6673, mul_34_17_n_6674, mul_34_17_n_6675,
     mul_34_17_n_6676, mul_34_17_n_6677, mul_34_17_n_6678, mul_34_17_n_6679,
     mul_34_17_n_6680, mul_34_17_n_6681, mul_34_17_n_6682, mul_34_17_n_6683,
     mul_34_17_n_6684, mul_34_17_n_6685, mul_34_17_n_6686, mul_34_17_n_6687,
     mul_34_17_n_6688, mul_34_17_n_6689, mul_34_17_n_6690, mul_34_17_n_6691,
     mul_34_17_n_6692, mul_34_17_n_6693, mul_34_17_n_6694, mul_34_17_n_6695,
     mul_34_17_n_6696, mul_34_17_n_6697, mul_34_17_n_6698, mul_34_17_n_6699,
     mul_34_17_n_6700, mul_34_17_n_6701, mul_34_17_n_6702, mul_34_17_n_6703,
     mul_34_17_n_6704, mul_34_17_n_6705, mul_34_17_n_6706, mul_34_17_n_6707,
     mul_34_17_n_6708, mul_34_17_n_6709, mul_34_17_n_6710, mul_34_17_n_6711,
     mul_34_17_n_6712, mul_34_17_n_6713, mul_34_17_n_6714, mul_34_17_n_6715,
     mul_34_17_n_6716, mul_34_17_n_6717, mul_34_17_n_6718, mul_34_17_n_6719,
     mul_34_17_n_6720, mul_34_17_n_6721, mul_34_17_n_6722, mul_34_17_n_6723,
     mul_34_17_n_6724, mul_34_17_n_6725, mul_34_17_n_6726, mul_34_17_n_6727,
     mul_34_17_n_6728, mul_34_17_n_6729, mul_34_17_n_6730, mul_34_17_n_6731,
     mul_34_17_n_6732, mul_34_17_n_6733, mul_34_17_n_6734, mul_34_17_n_6735,
     mul_34_17_n_6736, mul_34_17_n_6737, mul_34_17_n_6738, mul_34_17_n_6739,
     mul_34_17_n_6740, mul_34_17_n_6741, mul_34_17_n_6742, mul_34_17_n_6743,
     mul_34_17_n_6744, mul_34_17_n_6745, mul_34_17_n_6746, mul_34_17_n_6747,
     mul_34_17_n_6748, mul_34_17_n_6749, mul_34_17_n_6750, mul_34_17_n_6751,
     mul_34_17_n_6752, mul_34_17_n_6753, mul_34_17_n_6754, mul_34_17_n_6755,
     mul_34_17_n_6756, mul_34_17_n_6757, mul_34_17_n_6758, mul_34_17_n_6759,
     mul_34_17_n_6760, mul_34_17_n_6761, mul_34_17_n_6762, mul_34_17_n_6763,
     mul_34_17_n_6764, mul_34_17_n_6767, mul_34_17_n_6776, mul_34_17_n_6777,
     mul_34_17_n_6778, mul_34_17_n_6779, mul_34_17_n_6780, mul_34_17_n_6781,
     mul_34_17_n_6782, mul_34_17_n_6783, mul_34_17_n_6784, mul_34_17_n_6785,
     mul_34_17_n_6786, mul_34_17_n_6787, mul_34_17_n_6788, mul_34_17_n_6789,
     mul_34_17_n_6790, mul_34_17_n_6791, mul_34_17_n_6792, mul_34_17_n_6793,
     mul_34_17_n_6794, mul_34_17_n_6795, mul_34_17_n_6796, mul_34_17_n_6797,
     mul_34_17_n_6798, mul_34_17_n_6800, mul_34_17_n_6801, mul_34_17_n_6802,
     mul_34_17_n_6803, mul_34_17_n_6804, mul_34_17_n_6805, mul_34_17_n_6806,
     mul_34_17_n_6807, mul_34_17_n_6808, mul_34_17_n_6809, mul_34_17_n_6810,
     mul_34_17_n_6811, mul_34_17_n_6812, mul_34_17_n_6813, mul_34_17_n_6814,
     mul_34_17_n_6815, mul_34_17_n_6816, mul_34_17_n_6817, mul_34_17_n_6818,
     mul_34_17_n_6819, mul_34_17_n_6820, mul_34_17_n_6821, mul_34_17_n_6822,
     mul_34_17_n_6823, mul_34_17_n_6824, mul_34_17_n_6825, mul_34_17_n_6826,
     mul_34_17_n_6827, mul_34_17_n_6828, mul_34_17_n_6829, mul_34_17_n_6830,
     mul_34_17_n_6831, mul_34_17_n_6832, mul_34_17_n_6834, mul_34_17_n_6835,
     mul_34_17_n_6836, mul_34_17_n_6837, mul_34_17_n_6838, mul_34_17_n_6839,
     mul_34_17_n_6840, mul_34_17_n_6841, mul_34_17_n_6842, mul_34_17_n_6843,
     mul_34_17_n_6844, mul_34_17_n_6845, mul_34_17_n_6846, mul_34_17_n_6847,
     mul_34_17_n_6848, mul_34_17_n_6849, mul_34_17_n_6850, mul_34_17_n_6851,
     mul_34_17_n_6852, mul_34_17_n_6853, mul_34_17_n_6854, mul_34_17_n_6855,
     mul_34_17_n_6856, mul_34_17_n_6857, mul_34_17_n_6858, mul_34_17_n_6859,
     mul_34_17_n_6860, mul_34_17_n_6861, mul_34_17_n_6862, mul_34_17_n_6864,
     mul_34_17_n_6867, mul_34_17_n_6870, mul_34_17_n_6871, mul_34_17_n_6872,
     mul_34_17_n_6875, mul_34_17_n_6876, mul_34_17_n_6882, mul_34_17_n_6883,
     mul_34_17_n_6884, mul_34_17_n_6885, mul_34_17_n_6886, mul_34_17_n_6887,
     mul_34_17_n_6888, mul_34_17_n_6890, mul_34_17_n_6891, mul_34_17_n_6893,
     mul_34_17_n_6894, mul_34_17_n_6895, mul_34_17_n_6896, mul_34_17_n_6897,
     mul_34_17_n_6898, mul_34_17_n_6899, mul_34_17_n_6900, mul_34_17_n_6901,
     mul_34_17_n_6902, mul_34_17_n_6903, mul_34_17_n_6904, mul_34_17_n_6905,
     mul_34_17_n_6906, mul_34_17_n_6907, mul_34_17_n_6908, mul_34_17_n_6909,
     mul_34_17_n_6910, mul_34_17_n_6911, mul_34_17_n_6912, mul_34_17_n_6913,
     mul_34_17_n_6914, mul_34_17_n_6915, mul_34_17_n_6916, mul_34_17_n_6917,
     mul_34_17_n_6918, mul_34_17_n_6919, mul_34_17_n_6920, mul_34_17_n_6921,
     mul_34_17_n_6922, mul_34_17_n_6923, mul_34_17_n_6924, mul_34_17_n_6925,
     mul_34_17_n_6926, mul_34_17_n_6927, mul_34_17_n_6928, mul_34_17_n_6929,
     mul_34_17_n_6930, mul_34_17_n_6931, mul_34_17_n_6932, mul_34_17_n_6933,
     mul_34_17_n_6934, mul_34_17_n_6935, mul_34_17_n_6936, mul_34_17_n_6937,
     mul_34_17_n_6938, mul_34_17_n_6939, mul_34_17_n_6940, mul_34_17_n_6941,
     mul_34_17_n_6942, mul_34_17_n_6943, mul_34_17_n_6944, mul_34_17_n_6945,
     mul_34_17_n_6946, mul_34_17_n_6947, mul_34_17_n_6948, mul_34_17_n_6949,
     mul_34_17_n_6950, mul_34_17_n_6951, mul_34_17_n_6952, mul_34_17_n_6953,
     mul_34_17_n_6954, mul_34_17_n_6955, mul_34_17_n_6956, mul_34_17_n_6957,
     mul_34_17_n_6958, mul_34_17_n_6959, mul_34_17_n_6960, mul_34_17_n_6961,
     mul_34_17_n_6962, mul_34_17_n_6963, mul_34_17_n_6964, mul_34_17_n_6965,
     mul_34_17_n_6966, mul_34_17_n_6967, mul_34_17_n_6969, mul_34_17_n_6970,
     mul_34_17_n_6971, mul_34_17_n_6974, mul_34_17_n_6975, mul_34_17_n_6976,
     mul_34_17_n_6978, mul_34_17_n_6979, mul_34_17_n_6983, mul_34_17_n_6984,
     mul_34_17_n_6985, mul_34_17_n_6987, mul_34_17_n_6989, mul_34_17_n_6990,
     mul_34_17_n_6992, mul_34_17_n_6993, mul_34_17_n_6994, mul_34_17_n_6995,
     mul_34_17_n_7000, mul_34_17_n_7002, mul_34_17_n_7011, mul_34_17_n_7012,
     mul_34_17_n_7014, mul_34_17_n_7019, mul_34_17_n_7020, mul_34_17_n_7022,
     mul_34_17_n_7024, mul_34_17_n_7027, mul_34_17_n_7028, mul_34_17_n_7038,
     mul_34_17_n_7043, mul_34_17_n_7044, mul_34_17_n_7046, mul_34_17_n_7048,
     mul_34_17_n_7049, mul_34_17_n_7050, mul_34_17_n_7051, mul_34_17_n_7052,
     mul_34_17_n_7053, mul_34_17_n_7054, mul_34_17_n_7055, mul_34_17_n_7056,
     mul_34_17_n_7057, mul_34_17_n_7058, mul_34_17_n_7059, mul_34_17_n_7060,
     mul_34_17_n_7061, mul_34_17_n_7062, mul_34_17_n_7063, mul_34_17_n_7064,
     mul_34_17_n_7065, mul_34_17_n_7066, mul_34_17_n_7067, mul_34_17_n_7068,
     mul_34_17_n_7069, mul_34_17_n_7070, mul_34_17_n_7071, mul_34_17_n_7072,
     mul_34_17_n_7073, mul_34_17_n_7074, mul_34_17_n_7075, mul_34_17_n_7076,
     mul_34_17_n_7077, mul_34_17_n_7078, mul_34_17_n_7079, mul_34_17_n_7080,
     mul_34_17_n_7081, mul_34_17_n_7082, mul_34_17_n_7083, mul_34_17_n_7084,
     mul_34_17_n_7085, mul_34_17_n_7086, mul_34_17_n_7087, mul_34_17_n_7088,
     mul_34_17_n_7089, mul_34_17_n_7090, mul_34_17_n_7091, mul_34_17_n_7092,
     mul_34_17_n_7093, mul_34_17_n_7094, mul_34_17_n_7095, mul_34_17_n_7096,
     mul_34_17_n_7097, mul_34_17_n_7098, mul_34_17_n_7099, mul_34_17_n_7100,
     mul_34_17_n_7101, mul_34_17_n_7102, mul_34_17_n_7103, mul_34_17_n_7104,
     mul_34_17_n_7105, mul_34_17_n_7106, mul_34_17_n_7107, mul_34_17_n_7108,
     mul_34_17_n_7109, mul_34_17_n_7110, mul_34_17_n_7111, mul_34_17_n_7112,
     mul_34_17_n_7113, mul_34_17_n_7114, mul_34_17_n_7115, mul_34_17_n_7116,
     mul_34_17_n_7117, mul_34_17_n_7118, mul_34_17_n_7119, mul_34_17_n_7120,
     mul_34_17_n_7121, mul_34_17_n_7122, mul_34_17_n_7123, mul_34_17_n_7124,
     mul_34_17_n_7125, mul_34_17_n_7126, mul_34_17_n_7127, mul_34_17_n_7128,
     mul_34_17_n_7129, mul_34_17_n_7130, mul_34_17_n_7131, mul_34_17_n_7132,
     mul_34_17_n_7133, mul_34_17_n_7134, mul_34_17_n_7135, mul_34_17_n_7136,
     mul_34_17_n_7137, mul_34_17_n_7138, mul_34_17_n_7139, mul_34_17_n_7140,
     mul_34_17_n_7141, mul_34_17_n_7142, mul_34_17_n_7143, mul_34_17_n_7144,
     mul_34_17_n_7145, mul_34_17_n_7146, mul_34_17_n_7147, mul_34_17_n_7148,
     mul_34_17_n_7149, mul_34_17_n_7150, mul_34_17_n_7151, mul_34_17_n_7152,
     mul_34_17_n_7153, mul_34_17_n_7154, mul_34_17_n_7155, mul_34_17_n_7156,
     mul_34_17_n_7157, mul_34_17_n_7158, mul_34_17_n_7159, mul_34_17_n_7160,
     mul_34_17_n_7161, mul_34_17_n_7162, mul_34_17_n_7163, mul_34_17_n_7164,
     mul_34_17_n_7165, mul_34_17_n_7166, mul_34_17_n_7167, mul_34_17_n_7168,
     mul_34_17_n_7169, mul_34_17_n_7170, mul_34_17_n_7171, mul_34_17_n_7172,
     mul_34_17_n_7173, mul_34_17_n_7174, mul_34_17_n_7175, mul_34_17_n_7176,
     mul_34_17_n_7177, mul_34_17_n_7178, mul_34_17_n_7179, mul_34_17_n_7180,
     mul_34_17_n_7181, mul_34_17_n_7182, mul_34_17_n_7183, mul_34_17_n_7184,
     mul_34_17_n_7185, mul_34_17_n_7186, mul_34_17_n_7187, mul_34_17_n_7188,
     mul_34_17_n_7189, mul_34_17_n_7190, mul_34_17_n_7191, mul_34_17_n_7193,
     mul_34_17_n_7194, mul_34_17_n_7195, mul_34_17_n_7198, mul_34_17_n_7199,
     mul_34_17_n_7205, mul_34_17_n_7207, mul_34_17_n_7208, mul_34_17_n_7209,
     mul_34_17_n_7210, mul_34_17_n_7216, mul_34_17_n_7217, mul_34_17_n_7218,
     mul_34_17_n_7219, mul_34_17_n_7220, mul_34_17_n_7230, mul_34_17_n_7233,
     mul_34_17_n_7237, mul_34_17_n_7238, mul_34_17_n_7240, mul_34_17_n_7242,
     mul_34_17_n_7244, mul_34_17_n_7245, mul_34_17_n_7246, mul_34_17_n_7247,
     mul_34_17_n_7248, mul_34_17_n_7249, mul_34_17_n_7250, mul_34_17_n_7251,
     mul_34_17_n_7252, mul_34_17_n_7253, mul_34_17_n_7255, mul_34_17_n_7256,
     mul_34_17_n_7258, mul_34_17_n_7259, mul_34_17_n_7260, mul_34_17_n_7261,
     mul_34_17_n_7263, mul_34_17_n_7265, mul_34_17_n_7266, mul_34_17_n_7267,
     mul_34_17_n_7268, mul_34_17_n_7273, mul_34_17_n_7274, mul_34_17_n_7276,
     mul_34_17_n_7277, mul_34_17_n_7278, mul_34_17_n_7280, mul_34_17_n_7281,
     mul_34_17_n_7282, mul_34_17_n_7283, mul_34_17_n_7284, mul_34_17_n_7285,
     mul_34_17_n_7286, mul_34_17_n_7287, mul_34_17_n_7288, mul_34_17_n_7289,
     mul_34_17_n_7290, mul_34_17_n_7291, mul_34_17_n_7292, mul_34_17_n_7293,
     mul_34_17_n_7294, mul_34_17_n_7295, mul_34_17_n_7296, mul_34_17_n_7297,
     mul_34_17_n_7298, mul_34_17_n_7299, mul_34_17_n_7300, mul_34_17_n_7301,
     mul_34_17_n_7302, mul_34_17_n_7303, mul_34_17_n_7304, mul_34_17_n_7305,
     mul_34_17_n_7306, mul_34_17_n_7307, mul_34_17_n_7308, mul_34_17_n_7309,
     mul_34_17_n_7310, mul_34_17_n_7311, mul_34_17_n_7312, mul_34_17_n_7313,
     mul_34_17_n_7314, mul_34_17_n_7315, mul_34_17_n_7316, mul_34_17_n_7317,
     mul_34_17_n_7318, mul_34_17_n_7319, mul_34_17_n_7320, mul_34_17_n_7321,
     mul_34_17_n_7322, mul_34_17_n_7323, mul_34_17_n_7324, mul_34_17_n_7325,
     mul_34_17_n_7326, mul_34_17_n_7327, mul_34_17_n_7328, mul_34_17_n_7329,
     mul_34_17_n_7330, mul_34_17_n_7331, mul_34_17_n_7332, mul_34_17_n_7333,
     mul_34_17_n_7334, mul_34_17_n_7335, mul_34_17_n_7336, mul_34_17_n_7337,
     mul_34_17_n_7338, mul_34_17_n_7339, mul_34_17_n_7340, mul_34_17_n_7341,
     mul_34_17_n_7342, mul_34_17_n_7343, mul_34_17_n_7344, mul_34_17_n_7345,
     mul_34_17_n_7346, mul_34_17_n_7347, mul_34_17_n_7348, mul_34_17_n_7349,
     mul_34_17_n_7350, mul_34_17_n_7351, mul_34_17_n_7352, mul_34_17_n_7353,
     mul_34_17_n_7354, mul_34_17_n_7355, mul_34_17_n_7356, mul_34_17_n_7357,
     mul_34_17_n_7358, mul_34_17_n_7359, mul_34_17_n_7360, mul_34_17_n_7361,
     mul_34_17_n_7362, mul_34_17_n_7363, mul_34_17_n_7364, mul_34_17_n_7365,
     mul_34_17_n_7366, mul_34_17_n_7367, mul_34_17_n_7368, mul_34_17_n_7369,
     mul_34_17_n_7370, mul_34_17_n_7371, mul_34_17_n_7372, mul_34_17_n_7373,
     mul_34_17_n_7374, mul_34_17_n_7375, mul_34_17_n_7376, mul_34_17_n_7377,
     mul_34_17_n_7378, mul_34_17_n_7379, mul_34_17_n_7380, mul_34_17_n_7381,
     mul_34_17_n_7382, mul_34_17_n_7383, mul_34_17_n_7384, mul_34_17_n_7385,
     mul_34_17_n_7386, mul_34_17_n_7387, mul_34_17_n_7388, mul_34_17_n_7389,
     mul_34_17_n_7390, mul_34_17_n_7391, mul_34_17_n_7392, mul_34_17_n_7393,
     mul_34_17_n_7394, mul_34_17_n_7395, mul_34_17_n_7396, mul_34_17_n_7397,
     mul_34_17_n_7399, mul_34_17_n_7400, mul_34_17_n_7401, mul_34_17_n_7402,
     mul_34_17_n_7403, mul_34_17_n_7404, mul_34_17_n_7405, mul_34_17_n_7407,
     mul_34_17_n_7408, mul_34_17_n_7410, mul_34_17_n_7411, mul_34_17_n_7412,
     mul_34_17_n_7413, mul_34_17_n_7414, mul_34_17_n_7415, mul_34_17_n_7416,
     mul_34_17_n_7418, mul_34_17_n_7420, mul_34_17_n_7421, mul_34_17_n_7422,
     mul_34_17_n_7423, mul_34_17_n_7424, mul_34_17_n_7425, mul_34_17_n_7427,
     mul_34_17_n_7428, mul_34_17_n_7429, mul_34_17_n_7430, mul_34_17_n_7431,
     mul_34_17_n_7433, mul_34_17_n_7434, mul_34_17_n_7435, mul_34_17_n_7436,
     mul_34_17_n_7437, mul_34_17_n_7438, mul_34_17_n_7439, mul_34_17_n_7440,
     mul_34_17_n_7441, mul_34_17_n_7442, mul_34_17_n_7443, mul_34_17_n_7444,
     mul_34_17_n_7445, mul_34_17_n_7446, mul_34_17_n_7447, mul_34_17_n_7448,
     mul_34_17_n_7449, mul_34_17_n_7450, mul_34_17_n_7451, mul_34_17_n_7452,
     mul_34_17_n_7453, mul_34_17_n_7454, mul_34_17_n_7455, mul_34_17_n_7456,
     mul_34_17_n_7457, mul_34_17_n_7458, mul_34_17_n_7459, mul_34_17_n_7460,
     mul_34_17_n_7461, mul_34_17_n_7462, mul_34_17_n_7463, mul_34_17_n_7464,
     mul_34_17_n_7465, mul_34_17_n_7466, mul_34_17_n_7467, mul_34_17_n_7468,
     mul_34_17_n_7469, mul_34_17_n_7470, mul_34_17_n_7471, mul_34_17_n_7472,
     mul_34_17_n_7473, mul_34_17_n_7474, mul_34_17_n_7475, mul_34_17_n_7476,
     mul_34_17_n_7478, mul_34_17_n_7479, mul_34_17_n_7480, mul_34_17_n_7481,
     mul_34_17_n_7482, mul_34_17_n_7483, mul_34_17_n_7484, mul_34_17_n_7486,
     mul_34_17_n_7487, mul_34_17_n_7488, mul_34_17_n_7489, mul_34_17_n_7490,
     mul_34_17_n_7491, mul_34_17_n_7492, mul_34_17_n_7493, mul_34_17_n_7494,
     mul_34_17_n_7495, mul_34_17_n_7496, mul_34_17_n_7497, mul_34_17_n_7498,
     mul_34_17_n_7499, mul_34_17_n_7500, mul_34_17_n_7501, mul_34_17_n_7503,
     mul_34_17_n_7504, mul_34_17_n_7505, mul_34_17_n_7506, mul_34_17_n_7507,
     mul_34_17_n_7508, mul_34_17_n_7509, mul_34_17_n_7511, mul_34_17_n_7512,
     mul_34_17_n_7513, mul_34_17_n_7514, mul_34_17_n_7515, mul_34_17_n_7516,
     mul_34_17_n_7517, mul_34_17_n_7518, mul_34_17_n_7519, mul_34_17_n_7520,
     mul_34_17_n_7521, mul_34_17_n_7522, mul_34_17_n_7523, mul_34_17_n_7524,
     mul_34_17_n_7525, mul_34_17_n_7526, mul_34_17_n_7527, mul_34_17_n_7528,
     mul_34_17_n_7529, mul_34_17_n_7530, mul_34_17_n_7531, mul_34_17_n_7532,
     mul_34_17_n_7533, mul_34_17_n_7534, mul_34_17_n_7535, mul_34_17_n_7536,
     mul_34_17_n_7537, mul_34_17_n_7538, mul_34_17_n_7539, mul_34_17_n_7540,
     mul_34_17_n_7541, mul_34_17_n_7542, mul_34_17_n_7544, mul_34_17_n_7545,
     mul_34_17_n_7546, mul_34_17_n_7547, mul_34_17_n_7548, mul_34_17_n_7549,
     mul_34_17_n_7550, mul_34_17_n_7551, mul_34_17_n_7552, mul_34_17_n_7553,
     mul_34_17_n_7554, mul_34_17_n_7555, mul_34_17_n_7556, mul_34_17_n_7557,
     mul_34_17_n_7558, mul_34_17_n_7559, mul_34_17_n_7560, mul_34_17_n_7561,
     mul_34_17_n_7562, mul_34_17_n_7563, mul_34_17_n_7564, mul_34_17_n_7565,
     mul_34_17_n_7566, mul_34_17_n_7567, mul_34_17_n_7568, mul_34_17_n_7570,
     mul_34_17_n_7572, mul_34_17_n_7573, mul_34_17_n_7576, mul_34_17_n_7577,
     mul_34_17_n_7579, mul_34_17_n_7580, mul_34_17_n_7581, mul_34_17_n_7582,
     mul_34_17_n_7583, mul_34_17_n_7584, mul_34_17_n_7585, mul_34_17_n_7586,
     mul_34_17_n_7587, mul_34_17_n_7588, mul_34_17_n_7589, mul_34_17_n_7590,
     mul_34_17_n_7591, mul_34_17_n_7592, mul_34_17_n_7593, mul_34_17_n_7594,
     mul_34_17_n_7595, mul_34_17_n_7596, mul_34_17_n_7597, mul_34_17_n_7598,
     mul_34_17_n_7599, mul_34_17_n_7600, mul_34_17_n_7601, mul_34_17_n_7602,
     mul_34_17_n_7603, mul_34_17_n_7604, mul_34_17_n_7605, mul_34_17_n_7606,
     mul_34_17_n_7607, mul_34_17_n_7608, mul_34_17_n_7609, mul_34_17_n_7610,
     mul_34_17_n_7611, mul_34_17_n_7612, mul_34_17_n_7613, mul_34_17_n_7614,
     mul_34_17_n_7615, mul_34_17_n_7616, mul_34_17_n_7617, mul_34_17_n_7618,
     mul_34_17_n_7619, mul_34_17_n_7620, mul_34_17_n_7621, mul_34_17_n_7622,
     mul_34_17_n_7623, mul_34_17_n_7624, mul_34_17_n_7625, mul_34_17_n_7626,
     mul_34_17_n_7627, mul_34_17_n_7628, mul_34_17_n_7629, mul_34_17_n_7630,
     mul_34_17_n_7631, mul_34_17_n_7632, mul_34_17_n_7633, mul_34_17_n_7634,
     mul_34_17_n_7635, mul_34_17_n_7636, mul_34_17_n_7637, mul_34_17_n_7638,
     mul_34_17_n_7639, mul_34_17_n_7640, mul_34_17_n_7641, mul_34_17_n_7642,
     mul_34_17_n_7643, mul_34_17_n_7644, mul_34_17_n_7645, mul_34_17_n_7646,
     mul_34_17_n_7647, mul_34_17_n_7648, mul_34_17_n_7649, mul_34_17_n_7650,
     mul_34_17_n_7651, mul_34_17_n_7652, mul_34_17_n_7653, mul_34_17_n_7654,
     mul_34_17_n_7655, mul_34_17_n_7656, mul_34_17_n_7657, mul_34_17_n_7658,
     mul_34_17_n_7659, mul_34_17_n_7660, mul_34_17_n_7661, mul_34_17_n_7662,
     mul_34_17_n_7663, mul_34_17_n_7664, mul_34_17_n_7665, mul_34_17_n_7666,
     mul_34_17_n_7667, mul_34_17_n_7668, mul_34_17_n_7669, mul_34_17_n_7670,
     mul_34_17_n_7671, mul_34_17_n_7672, mul_34_17_n_7673, mul_34_17_n_7674,
     mul_34_17_n_7675, mul_34_17_n_7677, mul_34_17_n_7678, mul_34_17_n_7679,
     mul_34_17_n_7680, mul_34_17_n_7681, mul_34_17_n_7682, mul_34_17_n_7684,
     mul_34_17_n_7685, mul_34_17_n_7686, mul_34_17_n_7687, mul_34_17_n_7688,
     mul_34_17_n_7689, mul_34_17_n_7690, mul_34_17_n_7691, mul_34_17_n_7692,
     mul_34_17_n_7693, mul_34_17_n_7694, mul_34_17_n_7695, mul_34_17_n_7696,
     mul_34_17_n_7697, mul_34_17_n_7698, mul_34_17_n_7699, mul_34_17_n_7700,
     mul_34_17_n_7701, mul_34_17_n_7702, mul_34_17_n_7703, mul_34_17_n_7704,
     mul_34_17_n_7705, mul_34_17_n_7706, mul_34_17_n_7707, mul_34_17_n_7708,
     mul_34_17_n_7709, mul_34_17_n_7710, mul_34_17_n_7711, mul_34_17_n_7712,
     mul_34_17_n_7713, mul_34_17_n_7714, mul_34_17_n_7715, mul_34_17_n_7716,
     mul_34_17_n_7717, mul_34_17_n_7718, mul_34_17_n_7719, mul_34_17_n_7720,
     mul_34_17_n_7721, mul_34_17_n_7722, mul_34_17_n_7723, mul_34_17_n_7724,
     mul_34_17_n_7725, mul_34_17_n_7726, mul_34_17_n_7727, mul_34_17_n_7728,
     mul_34_17_n_7729, mul_34_17_n_7730, mul_34_17_n_7731, mul_34_17_n_7732,
     mul_34_17_n_7733, mul_34_17_n_7734, mul_34_17_n_7735, mul_34_17_n_7736,
     mul_34_17_n_7737, mul_34_17_n_7738, mul_34_17_n_7739, mul_34_17_n_7740,
     mul_34_17_n_7741, mul_34_17_n_7742, mul_34_17_n_7743, mul_34_17_n_7744,
     mul_34_17_n_7745, mul_34_17_n_7746, mul_34_17_n_7747, mul_34_17_n_7748,
     mul_34_17_n_7749, mul_34_17_n_7750, mul_34_17_n_7751, mul_34_17_n_7752,
     mul_34_17_n_7753, mul_34_17_n_7754, mul_34_17_n_7755, mul_34_17_n_7756,
     mul_34_17_n_7757, mul_34_17_n_7758, mul_34_17_n_7759, mul_34_17_n_7760,
     mul_34_17_n_7761, mul_34_17_n_7762, mul_34_17_n_7763, mul_34_17_n_7764,
     mul_34_17_n_7765, mul_34_17_n_7766, mul_34_17_n_7767, mul_34_17_n_7768,
     mul_34_17_n_7769, mul_34_17_n_7770, mul_34_17_n_7771, mul_34_17_n_7772,
     mul_34_17_n_7773, mul_34_17_n_7774, mul_34_17_n_7775, mul_34_17_n_7776,
     mul_34_17_n_7777, mul_34_17_n_7778, mul_34_17_n_7779, mul_34_17_n_7780,
     mul_34_17_n_7781, mul_34_17_n_7782, mul_34_17_n_7783, mul_34_17_n_7784,
     mul_34_17_n_7785, mul_34_17_n_7786, mul_34_17_n_7787, mul_34_17_n_7788,
     mul_34_17_n_7791, mul_34_17_n_7792, mul_34_17_n_7793, mul_34_17_n_7794,
     mul_34_17_n_7795, mul_34_17_n_7796, mul_34_17_n_7797, mul_34_17_n_7798,
     mul_34_17_n_7799, mul_34_17_n_7800, mul_34_17_n_7801, mul_34_17_n_7802,
     mul_34_17_n_7803, mul_34_17_n_7804, mul_34_17_n_7805, mul_34_17_n_7806,
     mul_34_17_n_7807, mul_34_17_n_7808, mul_34_17_n_7809, mul_34_17_n_7810,
     mul_34_17_n_7811, mul_34_17_n_7812, mul_34_17_n_7813, mul_34_17_n_7814,
     mul_34_17_n_7815, mul_34_17_n_7816, mul_34_17_n_7817, mul_34_17_n_7818,
     mul_34_17_n_7819, mul_34_17_n_7820, mul_34_17_n_7821, mul_34_17_n_7823,
     mul_34_17_n_7824, mul_34_17_n_7832, mul_34_17_n_7834, mul_34_17_n_7835,
     mul_34_17_n_7836, mul_34_17_n_7838, mul_34_17_n_7839, mul_34_17_n_7842,
     mul_34_17_n_7843, mul_34_17_n_7844, mul_34_17_n_7845, mul_34_17_n_7846,
     mul_34_17_n_7850, mul_34_17_n_7852, mul_34_17_n_7853, mul_34_17_n_7854,
     mul_34_17_n_7855, mul_34_17_n_7857, mul_34_17_n_7858, mul_34_17_n_7860,
     mul_34_17_n_7861, mul_34_17_n_7862, mul_34_17_n_7864, mul_34_17_n_7865,
     mul_34_17_n_7867, mul_34_17_n_7869, mul_34_17_n_7871, mul_34_17_n_7872,
     mul_34_17_n_7875, mul_34_17_n_7876, mul_34_17_n_7877, mul_34_17_n_7878,
     mul_34_17_n_7880, mul_34_17_n_7881, mul_34_17_n_7882, mul_34_17_n_7884,
     mul_34_17_n_7885, mul_34_17_n_7887, mul_34_17_n_7888, mul_34_17_n_7889,
     mul_34_17_n_7890, mul_34_17_n_7893, mul_34_17_n_7894, mul_34_17_n_7895,
     mul_34_17_n_7896, mul_34_17_n_7897, mul_34_17_n_7898, mul_34_17_n_7899,
     mul_34_17_n_7900, mul_34_17_n_7901, mul_34_17_n_7902, mul_34_17_n_7903,
     mul_34_17_n_7905, mul_34_17_n_7906, mul_34_17_n_7908, mul_34_17_n_7911,
     mul_34_17_n_7913, mul_34_17_n_7915, mul_34_17_n_7918, mul_34_17_n_7919,
     mul_34_17_n_7922, mul_34_17_n_7923, mul_34_17_n_7924, mul_34_17_n_7925,
     mul_34_17_n_7926, mul_34_17_n_7927, mul_34_17_n_7928, mul_34_17_n_7929,
     mul_34_17_n_7930, mul_34_17_n_7931, mul_34_17_n_7932, mul_34_17_n_7933,
     mul_34_17_n_7934, mul_34_17_n_7935, mul_34_17_n_7936, mul_34_17_n_7937,
     mul_34_17_n_7938, mul_34_17_n_7939, mul_34_17_n_7940, mul_34_17_n_7941,
     mul_34_17_n_7942, mul_34_17_n_7943, mul_34_17_n_7944, mul_34_17_n_7945,
     mul_34_17_n_7946, mul_34_17_n_7947, mul_34_17_n_7948, mul_34_17_n_7949,
     mul_34_17_n_7950, mul_34_17_n_7951, mul_34_17_n_7952, mul_34_17_n_7953,
     mul_34_17_n_7954, mul_34_17_n_7955, mul_34_17_n_7956, mul_34_17_n_7957,
     mul_34_17_n_7958, mul_34_17_n_7959, mul_34_17_n_7960, mul_34_17_n_7961,
     mul_34_17_n_7963, mul_34_17_n_7964, mul_34_17_n_7968, mul_34_17_n_7970,
     mul_34_17_n_7971, mul_34_17_n_7972, mul_34_17_n_7973, mul_34_17_n_7974,
     mul_34_17_n_7975, mul_34_17_n_7976, mul_34_17_n_7978, mul_34_17_n_7979,
     mul_34_17_n_7980, mul_34_17_n_7981, mul_34_17_n_7983, mul_34_17_n_7984,
     mul_34_17_n_7986, mul_34_17_n_7987, mul_34_17_n_7993, mul_34_17_n_7996,
     mul_34_17_n_7998, mul_34_17_n_8001, mul_34_17_n_8002, mul_34_17_n_8003,
     mul_34_17_n_8004, mul_34_17_n_8005, mul_34_17_n_8007, mul_34_17_n_8008,
     mul_34_17_n_8009, mul_34_17_n_8010, mul_34_17_n_8011, mul_34_17_n_8012,
     mul_34_17_n_8013, mul_34_17_n_8015, mul_34_17_n_8016, mul_34_17_n_8017,
     mul_34_17_n_8019, mul_34_17_n_8020, mul_34_17_n_8021, mul_34_17_n_8022,
     mul_34_17_n_8023, mul_34_17_n_8024, mul_34_17_n_8025, mul_34_17_n_8026,
     mul_34_17_n_8027, mul_34_17_n_8028, mul_34_17_n_8030, mul_34_17_n_8031,
     mul_34_17_n_8032, mul_34_17_n_8033, mul_34_17_n_8035, mul_34_17_n_8036,
     mul_34_17_n_8037, mul_34_17_n_8040, mul_34_17_n_8041, mul_34_17_n_8042,
     mul_34_17_n_8044, mul_34_17_n_8046, mul_34_17_n_8048, mul_34_17_n_8049,
     mul_34_17_n_8050, mul_34_17_n_8051, mul_34_17_n_8052, mul_34_17_n_8053,
     mul_34_17_n_8054, mul_34_17_n_8055, mul_34_17_n_8056, mul_34_17_n_8057,
     mul_34_17_n_8059, mul_34_17_n_8060, mul_34_17_n_8061, mul_34_17_n_8062,
     mul_34_17_n_8063, mul_34_17_n_8064, mul_34_17_n_8065, mul_34_17_n_8066,
     mul_34_17_n_8067, mul_34_17_n_8068, mul_34_17_n_8069, mul_34_17_n_8070,
     mul_34_17_n_8071, mul_34_17_n_8072, mul_34_17_n_8073, mul_34_17_n_8074,
     mul_34_17_n_8075, mul_34_17_n_8076, mul_34_17_n_8077, mul_34_17_n_8078,
     mul_34_17_n_8079, mul_34_17_n_8080, mul_34_17_n_8081, mul_34_17_n_8082,
     mul_34_17_n_8083, mul_34_17_n_8084, mul_34_17_n_8085, mul_34_17_n_8086,
     mul_34_17_n_8087, mul_34_17_n_8088, mul_34_17_n_8089, mul_34_17_n_8090,
     mul_34_17_n_8091, mul_34_17_n_8092, mul_34_17_n_8093, mul_34_17_n_8094,
     mul_34_17_n_8095, mul_34_17_n_8096, mul_34_17_n_8097, mul_34_17_n_8098,
     mul_34_17_n_8099, mul_34_17_n_8100, mul_34_17_n_8101, mul_34_17_n_8102,
     mul_34_17_n_8103, mul_34_17_n_8104, mul_34_17_n_8105, mul_34_17_n_8106,
     mul_34_17_n_8108, mul_34_17_n_8112, mul_34_17_n_8113, mul_34_17_n_8115,
     mul_34_17_n_8118, mul_34_17_n_8119, mul_34_17_n_8120, mul_34_17_n_8121,
     mul_34_17_n_8123, mul_34_17_n_8126, mul_34_17_n_8127, mul_34_17_n_8128,
     mul_34_17_n_8129, mul_34_17_n_8130, mul_34_17_n_8131, mul_34_17_n_8132,
     mul_34_17_n_8133, mul_34_17_n_8134, mul_34_17_n_8135, mul_34_17_n_8136,
     mul_34_17_n_8137, mul_34_17_n_8138, mul_34_17_n_8140, mul_34_17_n_8141,
     mul_34_17_n_8142, mul_34_17_n_8143, mul_34_17_n_8144, mul_34_17_n_8145,
     mul_34_17_n_8146, mul_34_17_n_8147, mul_34_17_n_8148, mul_34_17_n_8149,
     mul_34_17_n_8150, mul_34_17_n_8151, mul_34_17_n_8152, mul_34_17_n_8153,
     mul_34_17_n_8154, mul_34_17_n_8155, mul_34_17_n_8156, mul_34_17_n_8157,
     mul_34_17_n_8158, mul_34_17_n_8159, mul_34_17_n_8160, mul_34_17_n_8161,
     mul_34_17_n_8162, mul_34_17_n_8163, mul_34_17_n_8164, mul_34_17_n_8165,
     mul_34_17_n_8166, mul_34_17_n_8167, mul_34_17_n_8168, mul_34_17_n_8169,
     mul_34_17_n_8170, mul_34_17_n_8171, mul_34_17_n_8172, mul_34_17_n_8173,
     mul_34_17_n_8174, mul_34_17_n_8175, mul_34_17_n_8176, mul_34_17_n_8177,
     mul_34_17_n_8178, mul_34_17_n_8179, mul_34_17_n_8180, mul_34_17_n_8181,
     mul_34_17_n_8182, mul_34_17_n_8183, mul_34_17_n_8184, mul_34_17_n_8185,
     mul_34_17_n_8186, mul_34_17_n_8187, mul_34_17_n_8188, mul_34_17_n_8189,
     mul_34_17_n_8190, mul_34_17_n_8191, mul_34_17_n_8192, mul_34_17_n_8193,
     mul_34_17_n_8194, mul_34_17_n_8195, mul_34_17_n_8196, mul_34_17_n_8197,
     mul_34_17_n_8199, mul_34_17_n_8200, mul_34_17_n_8201, mul_34_17_n_8202,
     mul_34_17_n_8203, mul_34_17_n_8204, mul_34_17_n_8205, mul_34_17_n_8206,
     mul_34_17_n_8207, mul_34_17_n_8208, mul_34_17_n_8209, mul_34_17_n_8210,
     mul_34_17_n_8212, mul_34_17_n_8213, mul_34_17_n_8214, mul_34_17_n_8215,
     mul_34_17_n_8216, mul_34_17_n_8217, mul_34_17_n_8218, mul_34_17_n_8219,
     mul_34_17_n_8220, mul_34_17_n_8221, mul_34_17_n_8222, mul_34_17_n_8223,
     mul_34_17_n_8224, mul_34_17_n_8226, mul_34_17_n_8227, mul_34_17_n_8228,
     mul_34_17_n_8229, mul_34_17_n_8230, mul_34_17_n_8231, mul_34_17_n_8232,
     mul_34_17_n_8233, mul_34_17_n_8234, mul_34_17_n_8235, mul_34_17_n_8236,
     mul_34_17_n_8237, mul_34_17_n_8238, mul_34_17_n_8239, mul_34_17_n_8240,
     mul_34_17_n_8241, mul_34_17_n_8242, mul_34_17_n_8243, mul_34_17_n_8244,
     mul_34_17_n_8245, mul_34_17_n_8246, mul_34_17_n_8247, mul_34_17_n_8248,
     mul_34_17_n_8249, mul_34_17_n_8250, mul_34_17_n_8252, mul_34_17_n_8253,
     mul_34_17_n_8254, mul_34_17_n_8255, mul_34_17_n_8256, mul_34_17_n_8257,
     mul_34_17_n_8258, mul_34_17_n_8259, mul_34_17_n_8260, mul_34_17_n_8261,
     mul_34_17_n_8262, mul_34_17_n_8263, mul_34_17_n_8264, mul_34_17_n_8265,
     mul_34_17_n_8266, mul_34_17_n_8267, mul_34_17_n_8268, mul_34_17_n_8269,
     mul_34_17_n_8270, mul_34_17_n_8271, mul_34_17_n_8272, mul_34_17_n_8273,
     mul_34_17_n_8274, mul_34_17_n_8275, mul_34_17_n_8276, mul_34_17_n_8277,
     mul_34_17_n_8278, mul_34_17_n_8279, mul_34_17_n_8280, mul_34_17_n_8281,
     mul_34_17_n_8282, mul_34_17_n_8283, mul_34_17_n_8284, mul_34_17_n_8285,
     mul_34_17_n_8286, mul_34_17_n_8287, mul_34_17_n_8288, mul_34_17_n_8289,
     mul_34_17_n_8290, mul_34_17_n_8291, mul_34_17_n_8292, mul_34_17_n_8293,
     mul_34_17_n_8294, mul_34_17_n_8295, mul_34_17_n_8296, mul_34_17_n_8297,
     mul_34_17_n_8298, mul_34_17_n_8299, mul_34_17_n_8300, mul_34_17_n_8301,
     mul_34_17_n_8302, mul_34_17_n_8303, mul_34_17_n_8304, mul_34_17_n_8305,
     mul_34_17_n_8307, mul_34_17_n_8308, mul_34_17_n_8311, mul_34_17_n_8312,
     mul_34_17_n_8313, mul_34_17_n_8314, mul_34_17_n_8321, mul_34_17_n_8323,
     mul_34_17_n_8324, mul_34_17_n_8325, mul_34_17_n_8326, mul_34_17_n_8327,
     mul_34_17_n_8328, mul_34_17_n_8329, mul_34_17_n_8330, mul_34_17_n_8331,
     mul_34_17_n_8332, mul_34_17_n_8333, mul_34_17_n_8334, mul_34_17_n_8335,
     mul_34_17_n_8336, mul_34_17_n_8337, mul_34_17_n_8338, mul_34_17_n_8339,
     mul_34_17_n_8340, mul_34_17_n_8341, mul_34_17_n_8342, mul_34_17_n_8343,
     mul_34_17_n_8344, mul_34_17_n_8346, mul_34_17_n_8348, mul_34_17_n_8349,
     mul_34_17_n_8352, mul_34_17_n_8353, mul_34_17_n_8354, mul_34_17_n_8355,
     mul_34_17_n_8356, mul_34_17_n_8357, mul_34_17_n_8358, mul_34_17_n_8359,
     mul_34_17_n_8360, mul_34_17_n_8361, mul_34_17_n_8362, mul_34_17_n_8363,
     mul_34_17_n_8364, mul_34_17_n_8365, mul_34_17_n_8366, mul_34_17_n_8367,
     mul_34_17_n_8368, mul_34_17_n_8369, mul_34_17_n_8370, mul_34_17_n_8371,
     mul_34_17_n_8372, mul_34_17_n_8373, mul_34_17_n_8374, mul_34_17_n_8375,
     mul_34_17_n_8376, mul_34_17_n_8377, mul_34_17_n_8378, mul_34_17_n_8379,
     mul_34_17_n_8380, mul_34_17_n_8381, mul_34_17_n_8382, mul_34_17_n_8383,
     mul_34_17_n_8384, mul_34_17_n_8385, mul_34_17_n_8386, mul_34_17_n_8387,
     mul_34_17_n_8388, mul_34_17_n_8389, mul_34_17_n_8390, mul_34_17_n_8391,
     mul_34_17_n_8392, mul_34_17_n_8393, mul_34_17_n_8394, mul_34_17_n_8395,
     mul_34_17_n_8396, mul_34_17_n_8397, mul_34_17_n_8398, mul_34_17_n_8399,
     mul_34_17_n_8402, mul_34_17_n_8403, mul_34_17_n_8404, mul_34_17_n_8405,
     mul_34_17_n_8406, mul_34_17_n_8407, mul_34_17_n_8408, mul_34_17_n_8409,
     mul_34_17_n_8410, mul_34_17_n_8411, mul_34_17_n_8412, mul_34_17_n_8413,
     mul_34_17_n_8414, mul_34_17_n_8415, mul_34_17_n_8416, mul_34_17_n_8417,
     mul_34_17_n_8418, mul_34_17_n_8419, mul_34_17_n_8420, mul_34_17_n_8421,
     mul_34_17_n_8423, mul_34_17_n_8424, mul_34_17_n_8425, mul_34_17_n_8426,
     mul_34_17_n_8427, mul_34_17_n_8428, mul_34_17_n_8429, mul_34_17_n_8430,
     mul_34_17_n_8431, mul_34_17_n_8432, mul_34_17_n_8433, mul_34_17_n_8434,
     mul_34_17_n_8435, mul_34_17_n_8436, mul_34_17_n_8437, mul_34_17_n_8438,
     mul_34_17_n_8439, mul_34_17_n_8440, mul_34_17_n_8441, mul_34_17_n_8442,
     mul_34_17_n_8443, mul_34_17_n_8444, mul_34_17_n_8445, mul_34_17_n_8446,
     mul_34_17_n_8447, mul_34_17_n_8448, mul_34_17_n_8449, mul_34_17_n_8450,
     mul_34_17_n_8451, mul_34_17_n_8452, mul_34_17_n_8453, mul_34_17_n_8454,
     mul_34_17_n_8458, mul_34_17_n_8459, mul_34_17_n_8460, mul_34_17_n_8461,
     mul_34_17_n_8462, mul_34_17_n_8463, mul_34_17_n_8464, mul_34_17_n_8465,
     mul_34_17_n_8466, mul_34_17_n_8467, mul_34_17_n_8468, mul_34_17_n_8469,
     mul_34_17_n_8470, mul_34_17_n_8472, mul_34_17_n_8473, mul_34_17_n_8474,
     mul_34_17_n_8475, mul_34_17_n_8476, mul_34_17_n_8477, mul_34_17_n_8478,
     mul_34_17_n_8479, mul_34_17_n_8480, mul_34_17_n_8482, mul_34_17_n_8485,
     mul_34_17_n_8486, mul_34_17_n_8487, mul_34_17_n_8488, mul_34_17_n_8489,
     mul_34_17_n_8490, mul_34_17_n_8491, mul_34_17_n_8492, mul_34_17_n_8493,
     mul_34_17_n_8494, mul_34_17_n_8495, mul_34_17_n_8496, mul_34_17_n_8497,
     mul_34_17_n_8498, mul_34_17_n_8499, mul_34_17_n_8500, mul_34_17_n_8501,
     mul_34_17_n_8502, mul_34_17_n_8503, mul_34_17_n_8504, mul_34_17_n_8505,
     mul_34_17_n_8506, mul_34_17_n_8507, mul_34_17_n_8508, mul_34_17_n_8509,
     mul_34_17_n_8510, mul_34_17_n_8511, mul_34_17_n_8512, mul_34_17_n_8513,
     mul_34_17_n_8514, mul_34_17_n_8515, mul_34_17_n_8516, mul_34_17_n_8517,
     mul_34_17_n_8518, mul_34_17_n_8519, mul_34_17_n_8520, mul_34_17_n_8521,
     mul_34_17_n_8522, mul_34_17_n_8523, mul_34_17_n_8524, mul_34_17_n_8525,
     mul_34_17_n_8527, mul_34_17_n_8528, mul_34_17_n_8529, mul_34_17_n_8530,
     mul_34_17_n_8531, mul_34_17_n_8532, mul_34_17_n_8533, mul_34_17_n_8534,
     mul_34_17_n_8535, mul_34_17_n_8536, mul_34_17_n_8537, mul_34_17_n_8538,
     mul_34_17_n_8539, mul_34_17_n_8540, mul_34_17_n_8541, mul_34_17_n_8542,
     mul_34_17_n_8543, mul_34_17_n_8544, mul_34_17_n_8545, mul_34_17_n_8546,
     mul_34_17_n_8547, mul_34_17_n_8548, mul_34_17_n_8549, mul_34_17_n_8550,
     mul_34_17_n_8551, mul_34_17_n_8552, mul_34_17_n_8553, mul_34_17_n_8554,
     mul_34_17_n_8555, mul_34_17_n_8556, mul_34_17_n_8557, mul_34_17_n_8558,
     mul_34_17_n_8559, mul_34_17_n_8560, mul_34_17_n_8561, mul_34_17_n_8562,
     mul_34_17_n_8563, mul_34_17_n_8564, mul_34_17_n_8565, mul_34_17_n_8566,
     mul_34_17_n_8567, mul_34_17_n_8568, mul_34_17_n_8570, mul_34_17_n_8571,
     mul_34_17_n_8572, mul_34_17_n_8573, mul_34_17_n_8574, mul_34_17_n_8575,
     mul_34_17_n_8576, mul_34_17_n_8577, mul_34_17_n_8578, mul_34_17_n_8579,
     mul_34_17_n_8580, mul_34_17_n_8581, mul_34_17_n_8582, mul_34_17_n_8583,
     mul_34_17_n_8584, mul_34_17_n_8585, mul_34_17_n_8586, mul_34_17_n_8587,
     mul_34_17_n_8589, mul_34_17_n_8590, mul_34_17_n_8591, mul_34_17_n_8592,
     mul_34_17_n_8593, mul_34_17_n_8594, mul_34_17_n_8595, mul_34_17_n_8596,
     mul_34_17_n_8597, mul_34_17_n_8598, mul_34_17_n_8599, mul_34_17_n_8600,
     mul_34_17_n_8601, mul_34_17_n_8602, mul_34_17_n_8603, mul_34_17_n_8604,
     mul_34_17_n_8605, mul_34_17_n_8607, mul_34_17_n_8608, mul_34_17_n_8609,
     mul_34_17_n_8610, mul_34_17_n_8611, mul_34_17_n_8612, mul_34_17_n_8613,
     mul_34_17_n_8615, mul_34_17_n_8616, mul_34_17_n_8617, mul_34_17_n_8618,
     mul_34_17_n_8619, mul_34_17_n_8620, mul_34_17_n_8621, mul_34_17_n_8622,
     mul_34_17_n_8623, mul_34_17_n_8624, mul_34_17_n_8625, mul_34_17_n_8626,
     mul_34_17_n_8627, mul_34_17_n_8628, mul_34_17_n_8629, mul_34_17_n_8630,
     mul_34_17_n_8631, mul_34_17_n_8632, mul_34_17_n_8633, mul_34_17_n_8635,
     mul_34_17_n_8636, mul_34_17_n_8637, mul_34_17_n_8638, mul_34_17_n_8639,
     mul_34_17_n_8640, mul_34_17_n_8641, mul_34_17_n_8642, mul_34_17_n_8643,
     mul_34_17_n_8644, mul_34_17_n_8645, mul_34_17_n_8646, mul_34_17_n_8647,
     mul_34_17_n_8648, mul_34_17_n_8649, mul_34_17_n_8650, mul_34_17_n_8651,
     mul_34_17_n_8652, mul_34_17_n_8653, mul_34_17_n_8654, mul_34_17_n_8655,
     mul_34_17_n_8656, mul_34_17_n_8657, mul_34_17_n_8658, mul_34_17_n_8659,
     mul_34_17_n_8660, mul_34_17_n_8661, mul_34_17_n_8662, mul_34_17_n_8663,
     mul_34_17_n_8664, mul_34_17_n_8666, mul_34_17_n_8668, mul_34_17_n_8669,
     mul_34_17_n_8670, mul_34_17_n_8671, mul_34_17_n_8672, mul_34_17_n_8673,
     mul_34_17_n_8674, mul_34_17_n_8675, mul_34_17_n_8676, mul_34_17_n_8677,
     mul_34_17_n_8678, mul_34_17_n_8680, mul_34_17_n_8682, mul_34_17_n_8684,
     mul_34_17_n_8686, mul_34_17_n_8687, mul_34_17_n_8688, mul_34_17_n_8689,
     mul_34_17_n_8690, mul_34_17_n_8691, mul_34_17_n_8692, mul_34_17_n_8693,
     mul_34_17_n_8694, mul_34_17_n_8695, mul_34_17_n_8696, mul_34_17_n_8698,
     mul_34_17_n_8699, mul_34_17_n_8700, mul_34_17_n_8701, mul_34_17_n_8703,
     mul_34_17_n_8704, mul_34_17_n_8705, mul_34_17_n_8706, mul_34_17_n_8707,
     mul_34_17_n_8708, mul_34_17_n_8709, mul_34_17_n_8710, mul_34_17_n_8711,
     mul_34_17_n_8712, mul_34_17_n_8713, mul_34_17_n_8714, mul_34_17_n_8715,
     mul_34_17_n_8716, mul_34_17_n_8717, mul_34_17_n_8719, mul_34_17_n_8720,
     mul_34_17_n_8721, mul_34_17_n_8722, mul_34_17_n_8723, mul_34_17_n_8724,
     mul_34_17_n_8726, mul_34_17_n_8727, mul_34_17_n_8728, mul_34_17_n_8730,
     mul_34_17_n_8731, mul_34_17_n_8732, mul_34_17_n_8733, mul_34_17_n_8734,
     mul_34_17_n_8735, mul_34_17_n_8736, mul_34_17_n_8737, mul_34_17_n_8738,
     mul_34_17_n_8739, mul_34_17_n_8740, mul_34_17_n_8741, mul_34_17_n_8742,
     mul_34_17_n_8743, mul_34_17_n_8744, mul_34_17_n_8745, mul_34_17_n_8746,
     mul_34_17_n_8747, mul_34_17_n_8748, mul_34_17_n_8749, mul_34_17_n_8750,
     mul_34_17_n_8751, mul_34_17_n_8752, mul_34_17_n_8753, mul_34_17_n_8754,
     mul_34_17_n_8755, mul_34_17_n_8756, mul_34_17_n_8757, mul_34_17_n_8758,
     mul_34_17_n_8759, mul_34_17_n_8760, mul_34_17_n_8761, mul_34_17_n_8762,
     mul_34_17_n_8763, mul_34_17_n_8764, mul_34_17_n_8765, mul_34_17_n_8766,
     mul_34_17_n_8767, mul_34_17_n_8768, mul_34_17_n_8769, mul_34_17_n_8770,
     mul_34_17_n_8771, mul_34_17_n_8773, mul_34_17_n_8775, mul_34_17_n_8776,
     mul_34_17_n_8777, mul_34_17_n_8779, mul_34_17_n_8780, mul_34_17_n_8782,
     mul_34_17_n_8783, mul_34_17_n_8784, mul_34_17_n_8785, mul_34_17_n_8786,
     mul_34_17_n_8787, mul_34_17_n_8788, mul_34_17_n_8789, mul_34_17_n_8790,
     mul_34_17_n_8791, mul_34_17_n_8792, mul_34_17_n_8793, mul_34_17_n_8794,
     mul_34_17_n_8795, mul_34_17_n_8796, mul_34_17_n_8797, mul_34_17_n_8798,
     mul_34_17_n_8799, mul_34_17_n_8801, mul_34_17_n_8802, mul_34_17_n_8803,
     mul_34_17_n_8804, mul_34_17_n_8805, mul_34_17_n_8806, mul_34_17_n_8807,
     mul_34_17_n_8808, mul_34_17_n_8809, mul_34_17_n_8810, mul_34_17_n_8811,
     mul_34_17_n_8812, mul_34_17_n_8813, mul_34_17_n_8814, mul_34_17_n_8815,
     mul_34_17_n_8816, mul_34_17_n_8817, mul_34_17_n_8818, mul_34_17_n_8819,
     mul_34_17_n_8820, mul_34_17_n_8821, mul_34_17_n_8822, mul_34_17_n_8823,
     mul_34_17_n_8824, mul_34_17_n_8825, mul_34_17_n_8826, mul_34_17_n_8827,
     mul_34_17_n_8828, mul_34_17_n_8829, mul_34_17_n_8830, mul_34_17_n_8831,
     mul_34_17_n_8834, mul_34_17_n_8835, mul_34_17_n_8838, mul_34_17_n_8839,
     mul_34_17_n_8840, mul_34_17_n_8841, mul_34_17_n_8842, mul_34_17_n_8843,
     mul_34_17_n_8844, mul_34_17_n_8845, mul_34_17_n_8846, mul_34_17_n_8847,
     mul_34_17_n_8848, mul_34_17_n_8849, mul_34_17_n_8850, mul_34_17_n_8851,
     mul_34_17_n_8852, mul_34_17_n_8853, mul_34_17_n_8854, mul_34_17_n_8855,
     mul_34_17_n_8856, mul_34_17_n_8859, mul_34_17_n_8860, mul_34_17_n_8863,
     mul_34_17_n_8864, mul_34_17_n_8865, mul_34_17_n_8866, mul_34_17_n_8867,
     mul_34_17_n_8868, mul_34_17_n_8869, mul_34_17_n_8870, mul_34_17_n_8872,
     mul_34_17_n_8873, mul_34_17_n_8874, mul_34_17_n_8875, mul_34_17_n_8876,
     mul_34_17_n_8877, mul_34_17_n_8878, mul_34_17_n_8879, mul_34_17_n_8880,
     mul_34_17_n_8881, mul_34_17_n_8882, mul_34_17_n_8883, mul_34_17_n_8884,
     mul_34_17_n_8885, mul_34_17_n_8886, mul_34_17_n_8887, mul_34_17_n_8888,
     mul_34_17_n_8889, mul_34_17_n_8890, mul_34_17_n_8891, mul_34_17_n_8892,
     mul_34_17_n_8893, mul_34_17_n_8894, mul_34_17_n_8895, mul_34_17_n_8896,
     mul_34_17_n_8897, mul_34_17_n_8898, mul_34_17_n_8901, mul_34_17_n_8902,
     mul_34_17_n_8903, mul_34_17_n_8904, mul_34_17_n_8905, mul_34_17_n_8906,
     mul_34_17_n_8907, mul_34_17_n_8908, mul_34_17_n_8909, mul_34_17_n_8910,
     mul_34_17_n_8911, mul_34_17_n_8912, mul_34_17_n_8913, mul_34_17_n_8914,
     mul_34_17_n_8915, mul_34_17_n_8916, mul_34_17_n_8917, mul_34_17_n_8918,
     mul_34_17_n_8919, mul_34_17_n_8920, mul_34_17_n_8921, mul_34_17_n_8922,
     mul_34_17_n_8923, mul_34_17_n_8924, mul_34_17_n_8925, mul_34_17_n_8926,
     mul_34_17_n_8927, mul_34_17_n_8928, mul_34_17_n_8929, mul_34_17_n_8930,
     mul_34_17_n_8931, mul_34_17_n_8932, mul_34_17_n_8933, mul_34_17_n_8934,
     mul_34_17_n_8935, mul_34_17_n_8936, mul_34_17_n_8937, mul_34_17_n_8938,
     mul_34_17_n_8939, mul_34_17_n_8940, mul_34_17_n_8941, mul_34_17_n_8942,
     mul_34_17_n_8943, mul_34_17_n_8944, mul_34_17_n_8945, mul_34_17_n_8946,
     mul_34_17_n_8947, mul_34_17_n_8948, mul_34_17_n_8949, mul_34_17_n_8950,
     mul_34_17_n_8952, mul_34_17_n_8953, mul_34_17_n_8954, mul_34_17_n_8955,
     mul_34_17_n_8956, mul_34_17_n_8957, mul_34_17_n_8958, mul_34_17_n_8959,
     mul_34_17_n_8960, mul_34_17_n_8961, mul_34_17_n_8962, mul_34_17_n_8963,
     mul_34_17_n_8964, mul_34_17_n_8965, mul_34_17_n_8966, mul_34_17_n_8967,
     mul_34_17_n_8968, mul_34_17_n_8969, mul_34_17_n_8970, mul_34_17_n_8971,
     mul_34_17_n_8974, mul_34_17_n_8975, mul_34_17_n_8976, mul_34_17_n_8981,
     mul_34_17_n_8982, mul_34_17_n_8984, mul_34_17_n_8985, mul_34_17_n_8986,
     mul_34_17_n_8987, mul_34_17_n_8988, mul_34_17_n_8989, mul_34_17_n_8990,
     mul_34_17_n_8991, mul_34_17_n_8992, mul_34_17_n_8993, mul_34_17_n_8995,
     mul_34_17_n_8996, mul_34_17_n_8997, mul_34_17_n_8998, mul_34_17_n_8999,
     mul_34_17_n_9000, mul_34_17_n_9001, mul_34_17_n_9002, mul_34_17_n_9003,
     mul_34_17_n_9004, mul_34_17_n_9005, mul_34_17_n_9006, mul_34_17_n_9007,
     mul_34_17_n_9009, mul_34_17_n_9010, mul_34_17_n_9011, mul_34_17_n_9012,
     mul_34_17_n_9013, mul_34_17_n_9014, mul_34_17_n_9017, mul_34_17_n_9018,
     mul_34_17_n_9019, mul_34_17_n_9021, mul_34_17_n_9023, mul_34_17_n_9024,
     mul_34_17_n_9025, mul_34_17_n_9026, mul_34_17_n_9027, mul_34_17_n_9028,
     mul_34_17_n_9029, mul_34_17_n_9030, mul_34_17_n_9031, mul_34_17_n_9033,
     mul_34_17_n_9034, mul_34_17_n_9035, mul_34_17_n_9036, mul_34_17_n_9037,
     mul_34_17_n_9038, mul_34_17_n_9039, mul_34_17_n_9040, mul_34_17_n_9041,
     mul_34_17_n_9042, mul_34_17_n_9043, mul_34_17_n_9044, mul_34_17_n_9045,
     mul_34_17_n_9046, mul_34_17_n_9047, mul_34_17_n_9048, mul_34_17_n_9049,
     mul_34_17_n_9050, mul_34_17_n_9051, mul_34_17_n_9052, mul_34_17_n_9053,
     mul_34_17_n_9054, mul_34_17_n_9055, mul_34_17_n_9056, mul_34_17_n_9057,
     mul_34_17_n_9058, mul_34_17_n_9059, mul_34_17_n_9060, mul_34_17_n_9061,
     mul_34_17_n_9062, mul_34_17_n_9063, mul_34_17_n_9064, mul_34_17_n_9065,
     mul_34_17_n_9066, mul_34_17_n_9067, mul_34_17_n_9068, mul_34_17_n_9069,
     mul_34_17_n_9071, mul_34_17_n_9072, mul_34_17_n_9073, mul_34_17_n_9074,
     mul_34_17_n_9075, mul_34_17_n_9076, mul_34_17_n_9077, mul_34_17_n_9078,
     mul_34_17_n_9079, mul_34_17_n_9080, mul_34_17_n_9081, mul_34_17_n_9082,
     mul_34_17_n_9083, mul_34_17_n_9084, mul_34_17_n_9086, mul_34_17_n_9087,
     mul_34_17_n_9088, mul_34_17_n_9089, mul_34_17_n_9090, mul_34_17_n_9091,
     mul_34_17_n_9092, mul_34_17_n_9093, mul_34_17_n_9094, mul_34_17_n_9095,
     mul_34_17_n_9096, mul_34_17_n_9097, mul_34_17_n_9098, mul_34_17_n_9099,
     mul_34_17_n_9100, mul_34_17_n_9101, mul_34_17_n_9102, mul_34_17_n_9104,
     mul_34_17_n_9105, mul_34_17_n_9106, mul_34_17_n_9107, mul_34_17_n_9108,
     mul_34_17_n_9109, mul_34_17_n_9110, mul_34_17_n_9111, mul_34_17_n_9112,
     mul_34_17_n_9113, mul_34_17_n_9114, mul_34_17_n_9115, mul_34_17_n_9116,
     mul_34_17_n_9117, mul_34_17_n_9118, mul_34_17_n_9119, mul_34_17_n_9120,
     mul_34_17_n_9121, mul_34_17_n_9122, mul_34_17_n_9123, mul_34_17_n_9124,
     mul_34_17_n_9125, mul_34_17_n_9126, mul_34_17_n_9127, mul_34_17_n_9128,
     mul_34_17_n_9129, mul_34_17_n_9130, mul_34_17_n_9131, mul_34_17_n_9132,
     mul_34_17_n_9133, mul_34_17_n_9134, mul_34_17_n_9136, mul_34_17_n_9137,
     mul_34_17_n_9138, mul_34_17_n_9139, mul_34_17_n_9140, mul_34_17_n_9141,
     mul_34_17_n_9142, mul_34_17_n_9143, mul_34_17_n_9144, mul_34_17_n_9145,
     mul_34_17_n_9146, mul_34_17_n_9147, mul_34_17_n_9148, mul_34_17_n_9149,
     mul_34_17_n_9150, mul_34_17_n_9151, mul_34_17_n_9152, mul_34_17_n_9153,
     mul_34_17_n_9154, mul_34_17_n_9158, mul_34_17_n_9159, mul_34_17_n_9160,
     mul_34_17_n_9162, mul_34_17_n_9163, mul_34_17_n_9164, mul_34_17_n_9166,
     mul_34_17_n_9167, mul_34_17_n_9169, mul_34_17_n_9170, mul_34_17_n_9171,
     mul_34_17_n_9172, mul_34_17_n_9173, mul_34_17_n_9174, mul_34_17_n_9175,
     mul_34_17_n_9176, mul_34_17_n_9177, mul_34_17_n_9178, mul_34_17_n_9179,
     mul_34_17_n_9180, mul_34_17_n_9181, mul_34_17_n_9182, mul_34_17_n_9183,
     mul_34_17_n_9184, mul_34_17_n_9185, mul_34_17_n_9186, mul_34_17_n_9187,
     mul_34_17_n_9188, mul_34_17_n_9189, mul_34_17_n_9190, mul_34_17_n_9191,
     mul_34_17_n_9192, mul_34_17_n_9193, mul_34_17_n_9194, mul_34_17_n_9195,
     mul_34_17_n_9196, mul_34_17_n_9197, mul_34_17_n_9198, mul_34_17_n_9199,
     mul_34_17_n_9200, mul_34_17_n_9202, mul_34_17_n_9203, mul_34_17_n_9204,
     mul_34_17_n_9205, mul_34_17_n_9206, mul_34_17_n_9207, mul_34_17_n_9208,
     mul_34_17_n_9209, mul_34_17_n_9210, mul_34_17_n_9211, mul_34_17_n_9212,
     mul_34_17_n_9213, mul_34_17_n_9214, mul_34_17_n_9215, mul_34_17_n_9216,
     mul_34_17_n_9217, mul_34_17_n_9218, mul_34_17_n_9219, mul_34_17_n_9220,
     mul_34_17_n_9221, mul_34_17_n_9222, mul_34_17_n_9223, mul_34_17_n_9224,
     mul_34_17_n_9225, mul_34_17_n_9226, mul_34_17_n_9227, mul_34_17_n_9228,
     mul_34_17_n_9229, mul_34_17_n_9230, mul_34_17_n_9231, mul_34_17_n_9233,
     mul_34_17_n_9234, mul_34_17_n_9235, mul_34_17_n_9236, mul_34_17_n_9237,
     mul_34_17_n_9238, mul_34_17_n_9239, mul_34_17_n_9240, mul_34_17_n_9241,
     mul_34_17_n_9242, mul_34_17_n_9243, mul_34_17_n_9244, mul_34_17_n_9245,
     mul_34_17_n_9248, mul_34_17_n_9249, mul_34_17_n_9250, mul_34_17_n_9251,
     mul_34_17_n_9252, mul_34_17_n_9253, mul_34_17_n_9254, mul_34_17_n_9255,
     mul_34_17_n_9256, mul_34_17_n_9257, mul_34_17_n_9258, mul_34_17_n_9259,
     mul_34_17_n_9260, mul_34_17_n_9261, mul_34_17_n_9262, mul_34_17_n_9263,
     mul_34_17_n_9265, mul_34_17_n_9266, mul_34_17_n_9267, mul_34_17_n_9268,
     mul_34_17_n_9269, mul_34_17_n_9270, mul_34_17_n_9271, mul_34_17_n_9272,
     mul_34_17_n_9273, mul_34_17_n_9274, mul_34_17_n_9275, mul_34_17_n_9276,
     mul_34_17_n_9277, mul_34_17_n_9278, mul_34_17_n_9279, mul_34_17_n_9280,
     mul_34_17_n_9281, mul_34_17_n_9282, mul_34_17_n_9283, mul_34_17_n_9284,
     mul_34_17_n_9285, mul_34_17_n_9286, mul_34_17_n_9287, mul_34_17_n_9288,
     mul_34_17_n_9289, mul_34_17_n_9291, mul_34_17_n_9292, mul_34_17_n_9293,
     mul_34_17_n_9294, mul_34_17_n_9295, mul_34_17_n_9296, mul_34_17_n_9297,
     mul_34_17_n_9298, mul_34_17_n_9299, mul_34_17_n_9300, mul_34_17_n_9301,
     mul_34_17_n_9302, mul_34_17_n_9303, mul_34_17_n_9304, mul_34_17_n_9305,
     mul_34_17_n_9306, mul_34_17_n_9307, mul_34_17_n_9308, mul_34_17_n_9309,
     mul_34_17_n_9310, mul_34_17_n_9311, mul_34_17_n_9312, mul_34_17_n_9313,
     mul_34_17_n_9314, mul_34_17_n_9315, mul_34_17_n_9316, mul_34_17_n_9317,
     mul_34_17_n_9318, mul_34_17_n_9319, mul_34_17_n_9320, mul_34_17_n_9325,
     mul_34_17_n_9326, mul_34_17_n_9327, mul_34_17_n_9328, mul_34_17_n_9329,
     mul_34_17_n_9330, mul_34_17_n_9331, mul_34_17_n_9332, mul_34_17_n_9333,
     mul_34_17_n_9334, mul_34_17_n_9336, mul_34_17_n_9337, mul_34_17_n_9338,
     mul_34_17_n_9339, mul_34_17_n_9340, mul_34_17_n_9341, mul_34_17_n_9342,
     mul_34_17_n_9343, mul_34_17_n_9344, mul_34_17_n_9345, mul_34_17_n_9346,
     mul_34_17_n_9347, mul_34_17_n_9348, mul_34_17_n_9349, mul_34_17_n_9350,
     mul_34_17_n_9351, mul_34_17_n_9352, mul_34_17_n_9353, mul_34_17_n_9354,
     mul_34_17_n_9355, mul_34_17_n_9356, mul_34_17_n_9357, mul_34_17_n_9359,
     mul_34_17_n_9360, mul_34_17_n_9361, mul_34_17_n_9362, mul_34_17_n_9363,
     mul_34_17_n_9364, mul_34_17_n_9365, mul_34_17_n_9366, mul_34_17_n_9367,
     mul_34_17_n_9368, mul_34_17_n_9369, mul_34_17_n_9370, mul_34_17_n_9371,
     mul_34_17_n_9372, mul_34_17_n_9373, mul_34_17_n_9374, mul_34_17_n_9375,
     mul_34_17_n_9376, mul_34_17_n_9377, mul_34_17_n_9378, mul_34_17_n_9379,
     mul_34_17_n_9380, mul_34_17_n_9381, mul_34_17_n_9382, mul_34_17_n_9383,
     mul_34_17_n_9384, mul_34_17_n_9385, mul_34_17_n_9386, mul_34_17_n_9387,
     mul_34_17_n_9389, mul_34_17_n_9390, mul_34_17_n_9391, mul_34_17_n_9392,
     mul_34_17_n_9393, mul_34_17_n_9394, mul_34_17_n_9395, mul_34_17_n_9396,
     mul_34_17_n_9397, mul_34_17_n_9398, mul_34_17_n_9399, mul_34_17_n_9401,
     mul_34_17_n_9402, mul_34_17_n_9403, mul_34_17_n_9404, mul_34_17_n_9405,
     mul_34_17_n_9406, mul_34_17_n_9407, mul_34_17_n_9409, mul_34_17_n_9410,
     mul_34_17_n_9411, mul_34_17_n_9415, mul_34_17_n_9416, mul_34_17_n_9417,
     mul_34_17_n_9418, mul_34_17_n_9419, mul_34_17_n_9420, mul_34_17_n_9421,
     mul_34_17_n_9422, mul_34_17_n_9423, mul_34_17_n_9424, mul_34_17_n_9425,
     mul_34_17_n_9426, mul_34_17_n_9427, mul_34_17_n_9428, mul_34_17_n_9429,
     mul_34_17_n_9430, mul_34_17_n_9431, mul_34_17_n_9433, mul_34_17_n_9434,
     mul_34_17_n_9435, mul_34_17_n_9436, mul_34_17_n_9437, mul_34_17_n_9438,
     mul_34_17_n_9439, mul_34_17_n_9440, mul_34_17_n_9441, mul_34_17_n_9443,
     mul_34_17_n_9444, mul_34_17_n_9445, mul_34_17_n_9446, mul_34_17_n_9447,
     mul_34_17_n_9448, mul_34_17_n_9449, mul_34_17_n_9450, mul_34_17_n_9451,
     mul_34_17_n_9452, mul_34_17_n_9453, mul_34_17_n_9454, mul_34_17_n_9455,
     mul_34_17_n_9456, mul_34_17_n_9457, mul_34_17_n_9458, mul_34_17_n_9460,
     mul_34_17_n_9461, mul_34_17_n_9462, mul_34_17_n_9463, mul_34_17_n_9464,
     mul_34_17_n_9466, mul_34_17_n_9467, mul_34_17_n_9468, mul_34_17_n_9469,
     mul_34_17_n_9470, mul_34_17_n_9472, mul_34_17_n_9473, mul_34_17_n_9474,
     mul_34_17_n_9475, mul_34_17_n_9476, mul_34_17_n_9477, mul_34_17_n_9478,
     mul_34_17_n_9479, mul_34_17_n_9480, mul_34_17_n_9481, mul_34_17_n_9482,
     mul_34_17_n_9483, mul_34_17_n_9485, mul_34_17_n_9487, mul_34_17_n_9489,
     mul_34_17_n_9490, mul_34_17_n_9491, mul_34_17_n_9492, mul_34_17_n_9493,
     mul_34_17_n_9494, mul_34_17_n_9495, mul_34_17_n_9497, mul_34_17_n_9498,
     mul_34_17_n_9499, mul_34_17_n_9500, mul_34_17_n_9501, mul_34_17_n_9502,
     mul_34_17_n_9503, mul_34_17_n_9504, mul_34_17_n_9505, mul_34_17_n_9506,
     mul_34_17_n_9507, mul_34_17_n_9508, mul_34_17_n_9509, mul_34_17_n_9510,
     mul_34_17_n_9511, mul_34_17_n_9512, mul_34_17_n_9513, mul_34_17_n_9514,
     mul_34_17_n_9515, mul_34_17_n_9517, mul_34_17_n_9518, mul_34_17_n_9519,
     mul_34_17_n_9520, mul_34_17_n_9521, mul_34_17_n_9522, mul_34_17_n_9523,
     mul_34_17_n_9524, mul_34_17_n_9525, mul_34_17_n_9526, mul_34_17_n_9527,
     mul_34_17_n_9528, mul_34_17_n_9529, mul_34_17_n_9530, mul_34_17_n_9531,
     mul_34_17_n_9532, mul_34_17_n_9533, mul_34_17_n_9534, mul_34_17_n_9535,
     mul_34_17_n_9536, mul_34_17_n_9537, mul_34_17_n_9538, mul_34_17_n_9539,
     mul_34_17_n_9540, mul_34_17_n_9541, mul_34_17_n_9542, mul_34_17_n_9543,
     mul_34_17_n_9544, mul_34_17_n_9545, mul_34_17_n_9546, mul_34_17_n_9547,
     mul_34_17_n_9548, mul_34_17_n_9549, mul_34_17_n_9550, mul_34_17_n_9551,
     mul_34_17_n_9552, mul_34_17_n_9553, mul_34_17_n_9554, mul_34_17_n_9555,
     mul_34_17_n_9556, mul_34_17_n_9557, mul_34_17_n_9558, mul_34_17_n_9559,
     mul_34_17_n_9560, mul_34_17_n_9561, mul_34_17_n_9562, mul_34_17_n_9563,
     mul_34_17_n_9564, mul_34_17_n_9565, mul_34_17_n_9566, mul_34_17_n_9567,
     mul_34_17_n_9568, mul_34_17_n_9569, mul_34_17_n_9570, mul_34_17_n_9572,
     mul_34_17_n_9578, mul_34_17_n_9579, mul_34_17_n_9580, mul_34_17_n_9581,
     mul_34_17_n_9582, mul_34_17_n_9583, mul_34_17_n_9584, mul_34_17_n_9585,
     mul_34_17_n_9587, mul_34_17_n_9588, mul_34_17_n_9589, mul_34_17_n_9590,
     mul_34_17_n_9591, mul_34_17_n_9592, mul_34_17_n_9593, mul_34_17_n_9594,
     mul_34_17_n_9595, mul_34_17_n_9596, mul_34_17_n_9597, mul_34_17_n_9598,
     mul_34_17_n_9599, mul_34_17_n_9600, mul_34_17_n_9601, mul_34_17_n_9602,
     mul_34_17_n_9604, mul_34_17_n_9605, mul_34_17_n_9606, mul_34_17_n_9607,
     mul_34_17_n_9608, mul_34_17_n_9609, mul_34_17_n_9610, mul_34_17_n_9611,
     mul_34_17_n_9612, mul_34_17_n_9614, mul_34_17_n_9615, mul_34_17_n_9616,
     mul_34_17_n_9617, mul_34_17_n_9618, mul_34_17_n_9619, mul_34_17_n_9620,
     mul_34_17_n_9621, mul_34_17_n_9622, mul_34_17_n_9623, mul_34_17_n_9624,
     mul_34_17_n_9625, mul_34_17_n_9626, mul_34_17_n_9627, mul_34_17_n_9628,
     mul_34_17_n_9629, mul_34_17_n_9630, mul_34_17_n_9631, mul_34_17_n_9632,
     mul_34_17_n_9633, mul_34_17_n_9634, mul_34_17_n_9635, mul_34_17_n_9636,
     mul_34_17_n_9637, mul_34_17_n_9638, mul_34_17_n_9639, mul_34_17_n_9640,
     mul_34_17_n_9641, mul_34_17_n_9643, mul_34_17_n_9644, mul_34_17_n_9645,
     mul_34_17_n_9646, mul_34_17_n_9647, mul_34_17_n_9650, mul_34_17_n_9651,
     mul_34_17_n_9652, mul_34_17_n_9653, mul_34_17_n_9654, mul_34_17_n_9655,
     mul_34_17_n_9656, mul_34_17_n_9657, mul_34_17_n_9658, mul_34_17_n_9659,
     mul_34_17_n_9660, mul_34_17_n_9661, mul_34_17_n_9662, mul_34_17_n_9663,
     mul_34_17_n_9664, mul_34_17_n_9665, mul_34_17_n_9666, mul_34_17_n_9667,
     mul_34_17_n_9668, mul_34_17_n_9669, mul_34_17_n_9670, mul_34_17_n_9672,
     mul_34_17_n_9674, mul_34_17_n_9675, mul_34_17_n_9676, mul_34_17_n_9677,
     mul_34_17_n_9678, mul_34_17_n_9679, mul_34_17_n_9681, mul_34_17_n_9682,
     mul_34_17_n_9683, mul_34_17_n_9684, mul_34_17_n_9686, mul_34_17_n_9687,
     mul_34_17_n_9688, mul_34_17_n_9689, mul_34_17_n_9690, mul_34_17_n_9691,
     mul_34_17_n_9692, mul_34_17_n_9693, mul_34_17_n_9694, mul_34_17_n_9695,
     mul_34_17_n_9696, mul_34_17_n_9697, mul_34_17_n_9698, mul_34_17_n_9699,
     mul_34_17_n_9700, mul_34_17_n_9702, mul_34_17_n_9703, mul_34_17_n_9704,
     mul_34_17_n_9706, mul_34_17_n_9707, mul_34_17_n_9708, mul_34_17_n_9709,
     mul_34_17_n_9710, mul_34_17_n_9711, mul_34_17_n_9712, mul_34_17_n_9713,
     mul_34_17_n_9714, mul_34_17_n_9715, mul_34_17_n_9716, mul_34_17_n_9717,
     mul_34_17_n_9718, mul_34_17_n_9719, mul_34_17_n_9720, mul_34_17_n_9721,
     mul_34_17_n_9722, mul_34_17_n_9723, mul_34_17_n_9724, mul_34_17_n_9725,
     mul_34_17_n_9726, mul_34_17_n_9727, mul_34_17_n_9728, mul_34_17_n_9729,
     mul_34_17_n_9730, mul_34_17_n_9731, mul_34_17_n_9732, mul_34_17_n_9733,
     mul_34_17_n_9734, mul_34_17_n_9735, mul_34_17_n_9737, mul_34_17_n_9738,
     mul_34_17_n_9739, mul_34_17_n_9740, mul_34_17_n_9741, mul_34_17_n_9742,
     mul_34_17_n_9743, mul_34_17_n_9744, mul_34_17_n_9745, mul_34_17_n_9746,
     mul_34_17_n_9747, mul_34_17_n_9748, mul_34_17_n_9749, mul_34_17_n_9750,
     mul_34_17_n_9751, mul_34_17_n_9752, mul_34_17_n_9753, mul_34_17_n_9754,
     mul_34_17_n_9755, mul_34_17_n_9756, mul_34_17_n_9757, mul_34_17_n_9758,
     mul_34_17_n_9760, mul_34_17_n_9761, mul_34_17_n_9762, mul_34_17_n_9763,
     mul_34_17_n_9764, mul_34_17_n_9765, mul_34_17_n_9766, mul_34_17_n_9767,
     mul_34_17_n_9768, mul_34_17_n_9770, mul_34_17_n_9771, mul_34_17_n_9772,
     mul_34_17_n_9773, mul_34_17_n_9774, mul_34_17_n_9775, mul_34_17_n_9776,
     mul_34_17_n_9777, mul_34_17_n_9778, mul_34_17_n_9779, mul_34_17_n_9780,
     mul_34_17_n_9781, mul_34_17_n_9782, mul_34_17_n_9783, mul_34_17_n_9784,
     mul_34_17_n_9785, mul_34_17_n_9786, mul_34_17_n_9787, mul_34_17_n_9788,
     mul_34_17_n_9789, mul_34_17_n_9790, mul_34_17_n_9791, mul_34_17_n_9792,
     mul_34_17_n_9793, mul_34_17_n_9794, mul_34_17_n_9795, mul_34_17_n_9796,
     mul_34_17_n_9797, mul_34_17_n_9798, mul_34_17_n_9799, mul_34_17_n_9800,
     mul_34_17_n_9801, mul_34_17_n_9802, mul_34_17_n_9803, mul_34_17_n_9804,
     mul_34_17_n_9805, mul_34_17_n_9806, mul_34_17_n_9807, mul_34_17_n_9808,
     mul_34_17_n_9809, mul_34_17_n_9811, mul_34_17_n_9815, mul_34_17_n_9816,
     mul_34_17_n_9817, mul_34_17_n_9818, mul_34_17_n_9819, mul_34_17_n_9820,
     mul_34_17_n_9821, mul_34_17_n_9822, mul_34_17_n_9823, mul_34_17_n_9824,
     mul_34_17_n_9825, mul_34_17_n_9827, mul_34_17_n_9828, mul_34_17_n_9829,
     mul_34_17_n_9830, mul_34_17_n_9831, mul_34_17_n_9832, mul_34_17_n_9833,
     mul_34_17_n_9834, mul_34_17_n_9835, mul_34_17_n_9836, mul_34_17_n_9837,
     mul_34_17_n_9838, mul_34_17_n_9839, mul_34_17_n_9840, mul_34_17_n_9841,
     mul_34_17_n_9842, mul_34_17_n_9843, mul_34_17_n_9844, mul_34_17_n_9845,
     mul_34_17_n_9846, mul_34_17_n_9847, mul_34_17_n_9848, mul_34_17_n_9849,
     mul_34_17_n_9850, mul_34_17_n_9851, mul_34_17_n_9852, mul_34_17_n_9853,
     mul_34_17_n_9854, mul_34_17_n_9855, mul_34_17_n_9856, mul_34_17_n_9857,
     mul_34_17_n_9858, mul_34_17_n_9859, mul_34_17_n_9860, mul_34_17_n_9861,
     mul_34_17_n_9862, mul_34_17_n_9863, mul_34_17_n_9864, mul_34_17_n_9865,
     mul_34_17_n_9866, mul_34_17_n_9867, mul_34_17_n_9868, mul_34_17_n_9869,
     mul_34_17_n_9870, mul_34_17_n_9871, mul_34_17_n_9872, mul_34_17_n_9873,
     mul_34_17_n_9874, mul_34_17_n_9875, mul_34_17_n_9876, mul_34_17_n_9877,
     mul_34_17_n_9878, mul_34_17_n_9879, mul_34_17_n_9880, mul_34_17_n_9881,
     mul_34_17_n_9882, mul_34_17_n_9883, mul_34_17_n_9884, mul_34_17_n_9885,
     mul_34_17_n_9886, mul_34_17_n_9887, mul_34_17_n_9888, mul_34_17_n_9889,
     mul_34_17_n_9890, mul_34_17_n_9891, mul_34_17_n_9892, mul_34_17_n_9893,
     mul_34_17_n_9894, mul_34_17_n_9895, mul_34_17_n_9896, mul_34_17_n_9897,
     mul_34_17_n_9898, mul_34_17_n_9899, mul_34_17_n_9900, mul_34_17_n_9901,
     mul_34_17_n_9902, mul_34_17_n_9903, mul_34_17_n_9905, mul_34_17_n_9906,
     mul_34_17_n_9907, mul_34_17_n_9908, mul_34_17_n_9909, mul_34_17_n_9910,
     mul_34_17_n_9911, mul_34_17_n_9913, mul_34_17_n_9914, mul_34_17_n_9915,
     mul_34_17_n_9916, mul_34_17_n_9917, mul_34_17_n_9918, mul_34_17_n_9919,
     mul_34_17_n_9920, mul_34_17_n_9921, mul_34_17_n_9922, mul_34_17_n_9923,
     mul_34_17_n_9924, mul_34_17_n_9925, mul_34_17_n_9926, mul_34_17_n_9927,
     mul_34_17_n_9928, mul_34_17_n_9929, mul_34_17_n_9930, mul_34_17_n_9931,
     mul_34_17_n_9932, mul_34_17_n_9933, mul_34_17_n_9934, mul_34_17_n_9935,
     mul_34_17_n_9936, mul_34_17_n_9937, mul_34_17_n_9938, mul_34_17_n_9939,
     mul_34_17_n_9940, mul_34_17_n_9941, mul_34_17_n_9942, mul_34_17_n_9943,
     mul_34_17_n_9945, mul_34_17_n_9947, mul_34_17_n_9948, mul_34_17_n_9949,
     mul_34_17_n_9950, mul_34_17_n_9951, mul_34_17_n_9953, mul_34_17_n_9954,
     mul_34_17_n_9955, mul_34_17_n_9957, mul_34_17_n_9958, mul_34_17_n_9959,
     mul_34_17_n_9960, mul_34_17_n_9961, mul_34_17_n_9962, mul_34_17_n_9963,
     mul_34_17_n_9964, mul_34_17_n_9965, mul_34_17_n_9966, mul_34_17_n_9967,
     mul_34_17_n_9968, mul_34_17_n_9969, mul_34_17_n_9970, mul_34_17_n_9971,
     mul_34_17_n_9972, mul_34_17_n_9973, mul_34_17_n_9974, mul_34_17_n_9975,
     mul_34_17_n_9976, mul_34_17_n_9977, mul_34_17_n_9978, mul_34_17_n_9979,
     mul_34_17_n_9980, mul_34_17_n_9981, mul_34_17_n_9982, mul_34_17_n_9983,
     mul_34_17_n_9984, mul_34_17_n_9985, mul_34_17_n_9986, mul_34_17_n_9987,
     mul_34_17_n_9988, mul_34_17_n_9989, mul_34_17_n_9990, mul_34_17_n_9991,
     mul_34_17_n_9992, mul_34_17_n_9993, mul_34_17_n_9994, mul_34_17_n_9995,
     mul_34_17_n_9996, mul_34_17_n_9997, mul_34_17_n_9998, mul_34_17_n_9999,
     mul_34_17_n_10000, mul_34_17_n_10001, mul_34_17_n_10002, mul_34_17_n_10003,
     mul_34_17_n_10004, mul_34_17_n_10005, mul_34_17_n_10006, mul_34_17_n_10007,
     mul_34_17_n_10008, mul_34_17_n_10009, mul_34_17_n_10010, mul_34_17_n_10011,
     mul_34_17_n_10012, mul_34_17_n_10013, mul_34_17_n_10014, mul_34_17_n_10015,
     mul_34_17_n_10016, mul_34_17_n_10017, mul_34_17_n_10018, mul_34_17_n_10019,
     mul_34_17_n_10020, mul_34_17_n_10021, mul_34_17_n_10022, mul_34_17_n_10023,
     mul_34_17_n_10024, mul_34_17_n_10025, mul_34_17_n_10026, mul_34_17_n_10027,
     mul_34_17_n_10028, mul_34_17_n_10029, mul_34_17_n_10030, mul_34_17_n_10031,
     mul_34_17_n_10032, mul_34_17_n_10033, mul_34_17_n_10034, mul_34_17_n_10035,
     mul_34_17_n_10036, mul_34_17_n_10037, mul_34_17_n_10038, mul_34_17_n_10039,
     mul_34_17_n_10040, mul_34_17_n_10041, mul_34_17_n_10042, mul_34_17_n_10043,
     mul_34_17_n_10044, mul_34_17_n_10045, mul_34_17_n_10046, mul_34_17_n_10047,
     mul_34_17_n_10048, mul_34_17_n_10049, mul_34_17_n_10050, mul_34_17_n_10051,
     mul_34_17_n_10052, mul_34_17_n_10053, mul_34_17_n_10054, mul_34_17_n_10055,
     mul_34_17_n_10056, mul_34_17_n_10057, mul_34_17_n_10058, mul_34_17_n_10059,
     mul_34_17_n_10060, mul_34_17_n_10061, mul_34_17_n_10062, mul_34_17_n_10063,
     mul_34_17_n_10064, mul_34_17_n_10065, mul_34_17_n_10066, mul_34_17_n_10067,
     mul_34_17_n_10068, mul_34_17_n_10069, mul_34_17_n_10071, mul_34_17_n_10072,
     mul_34_17_n_10073, mul_34_17_n_10074, mul_34_17_n_10075, mul_34_17_n_10076,
     mul_34_17_n_10077, mul_34_17_n_10078, mul_34_17_n_10079, mul_34_17_n_10080,
     mul_34_17_n_10081, mul_34_17_n_10082, mul_34_17_n_10083, mul_34_17_n_10084,
     mul_34_17_n_10085, mul_34_17_n_10086, mul_34_17_n_10087, mul_34_17_n_10088,
     mul_34_17_n_10089, mul_34_17_n_10090, mul_34_17_n_10091, mul_34_17_n_10092,
     mul_34_17_n_10093, mul_34_17_n_10094, mul_34_17_n_10095, mul_34_17_n_10096,
     mul_34_17_n_10097, mul_34_17_n_10098, mul_34_17_n_10099, mul_34_17_n_10100,
     mul_34_17_n_10101, mul_34_17_n_10102, mul_34_17_n_10103, mul_34_17_n_10104,
     mul_34_17_n_10105, mul_34_17_n_10106, mul_34_17_n_10107, mul_34_17_n_10108,
     mul_34_17_n_10109, mul_34_17_n_10110, mul_34_17_n_10111, mul_34_17_n_10112,
     mul_34_17_n_10113, mul_34_17_n_10114, mul_34_17_n_10115, mul_34_17_n_10116,
     mul_34_17_n_10117, mul_34_17_n_10118, mul_34_17_n_10119, mul_34_17_n_10120,
     mul_34_17_n_10121, mul_34_17_n_10122, mul_34_17_n_10123, mul_34_17_n_10124,
     mul_34_17_n_10125, mul_34_17_n_10126, mul_34_17_n_10127, mul_34_17_n_10128,
     mul_34_17_n_10129, mul_34_17_n_10130, mul_34_17_n_10131, mul_34_17_n_10132,
     mul_34_17_n_10133, mul_34_17_n_10134, mul_34_17_n_10135, mul_34_17_n_10136,
     mul_34_17_n_10137, mul_34_17_n_10138, mul_34_17_n_10139, mul_34_17_n_10140,
     mul_34_17_n_10141, mul_34_17_n_10142, mul_34_17_n_10143, mul_34_17_n_10144,
     mul_34_17_n_10145, mul_34_17_n_10146, mul_34_17_n_10147, mul_34_17_n_10148,
     mul_34_17_n_10149, mul_34_17_n_10150, mul_34_17_n_10151, mul_34_17_n_10152,
     mul_34_17_n_10153, mul_34_17_n_10154, mul_34_17_n_10155, mul_34_17_n_10156,
     mul_34_17_n_10157, mul_34_17_n_10158, mul_34_17_n_10159, mul_34_17_n_10160,
     mul_34_17_n_10161, mul_34_17_n_10162, mul_34_17_n_10163, mul_34_17_n_10164,
     mul_34_17_n_10165, mul_34_17_n_10166, mul_34_17_n_10167, mul_34_17_n_10168,
     mul_34_17_n_10169, mul_34_17_n_10170, mul_34_17_n_10171, mul_34_17_n_10172,
     mul_34_17_n_10173, mul_34_17_n_10174, mul_34_17_n_10175, mul_34_17_n_10176,
     mul_34_17_n_10177, mul_34_17_n_10178, mul_34_17_n_10179, mul_34_17_n_10180,
     mul_34_17_n_10181, mul_34_17_n_10182, mul_34_17_n_10183, mul_34_17_n_10184,
     mul_34_17_n_10185, mul_34_17_n_10186, mul_34_17_n_10187, mul_34_17_n_10188,
     mul_34_17_n_10189, mul_34_17_n_10190, mul_34_17_n_10191, mul_34_17_n_10192,
     mul_34_17_n_10193, mul_34_17_n_10194, mul_34_17_n_10195, mul_34_17_n_10196,
     mul_34_17_n_10197, mul_34_17_n_10198, mul_34_17_n_10199, mul_34_17_n_10200,
     mul_34_17_n_10201, mul_34_17_n_10202, mul_34_17_n_10203, mul_34_17_n_10204,
     mul_34_17_n_10205, mul_34_17_n_10206, mul_34_17_n_10207, mul_34_17_n_10208,
     mul_34_17_n_10209, mul_34_17_n_10210, mul_34_17_n_10211, mul_34_17_n_10212,
     mul_34_17_n_10213, mul_34_17_n_10214, mul_34_17_n_10215, mul_34_17_n_10216,
     mul_34_17_n_10217, mul_34_17_n_10218, mul_34_17_n_10219, mul_34_17_n_10220,
     mul_34_17_n_10221, mul_34_17_n_10222, mul_34_17_n_10223, mul_34_17_n_10224,
     mul_34_17_n_10225, mul_34_17_n_10226, mul_34_17_n_10227, mul_34_17_n_10228,
     mul_34_17_n_10229, mul_34_17_n_10230, mul_34_17_n_10231, mul_34_17_n_10232,
     mul_34_17_n_10233, mul_34_17_n_10234, mul_34_17_n_10235, mul_34_17_n_10236,
     mul_34_17_n_10237, mul_34_17_n_10238, mul_34_17_n_10239, mul_34_17_n_10240,
     mul_34_17_n_10241, mul_34_17_n_10242, mul_34_17_n_10243, mul_34_17_n_10244,
     mul_34_17_n_10245, mul_34_17_n_10246, mul_34_17_n_10247, mul_34_17_n_10248,
     mul_34_17_n_10249, mul_34_17_n_10250, mul_34_17_n_10251, mul_34_17_n_10252,
     mul_34_17_n_10253, mul_34_17_n_10254, mul_34_17_n_10255, mul_34_17_n_10256,
     mul_34_17_n_10257, mul_34_17_n_10258, mul_34_17_n_10259, mul_34_17_n_10260,
     mul_34_17_n_10261, mul_34_17_n_10262, mul_34_17_n_10263, mul_34_17_n_10264,
     mul_34_17_n_10265, mul_34_17_n_10266, mul_34_17_n_10267, mul_34_17_n_10268,
     mul_34_17_n_10269, mul_34_17_n_10270, mul_34_17_n_10271, mul_34_17_n_10272,
     mul_34_17_n_10273, mul_34_17_n_10274, mul_34_17_n_10275, mul_34_17_n_10276,
     mul_34_17_n_10277, mul_34_17_n_10278, mul_34_17_n_10279, mul_34_17_n_10280,
     mul_34_17_n_10281, mul_34_17_n_10282, mul_34_17_n_10283, mul_34_17_n_10284,
     mul_34_17_n_10285, mul_34_17_n_10286, mul_34_17_n_10287, mul_34_17_n_10288,
     mul_34_17_n_10289, mul_34_17_n_10290, mul_34_17_n_10291, mul_34_17_n_10292,
     mul_34_17_n_10293, mul_34_17_n_10294, mul_34_17_n_10295, mul_34_17_n_10296,
     mul_34_17_n_10297, mul_34_17_n_10298, mul_34_17_n_10299, mul_34_17_n_10300,
     mul_34_17_n_10301, mul_34_17_n_10302, mul_34_17_n_10303, mul_34_17_n_10304,
     mul_34_17_n_10305, mul_34_17_n_10306, mul_34_17_n_10307, mul_34_17_n_10308,
     mul_34_17_n_10309, mul_34_17_n_10310, mul_34_17_n_10311, mul_34_17_n_10312,
     mul_34_17_n_10313, mul_34_17_n_10314, mul_34_17_n_10315, mul_34_17_n_10316,
     mul_34_17_n_10317, mul_34_17_n_10318, mul_34_17_n_10319, mul_34_17_n_10320,
     mul_34_17_n_10321, mul_34_17_n_10322, mul_34_17_n_10323, mul_34_17_n_10324,
     mul_34_17_n_10325, mul_34_17_n_10326, mul_34_17_n_10327, mul_34_17_n_10328,
     mul_34_17_n_10329, mul_34_17_n_10330, mul_34_17_n_10331, mul_34_17_n_10332,
     mul_34_17_n_10333, mul_34_17_n_10334, mul_34_17_n_10335, mul_34_17_n_10336,
     mul_34_17_n_10337, mul_34_17_n_10338, mul_34_17_n_10339, mul_34_17_n_10340,
     mul_34_17_n_10341, mul_34_17_n_10342, mul_34_17_n_10343, mul_34_17_n_10344,
     mul_34_17_n_10345, mul_34_17_n_10346, mul_34_17_n_10347, mul_34_17_n_10348,
     mul_34_17_n_10349, mul_34_17_n_10350, mul_34_17_n_10351, mul_34_17_n_10352,
     mul_34_17_n_10353, mul_34_17_n_10354, mul_34_17_n_10355, mul_34_17_n_10356,
     mul_34_17_n_10357, mul_34_17_n_10358, mul_34_17_n_10359, mul_34_17_n_10360,
     mul_34_17_n_10361, mul_34_17_n_10362, mul_34_17_n_10363, mul_34_17_n_10364,
     mul_34_17_n_10365, mul_34_17_n_10366, mul_34_17_n_10367, mul_34_17_n_10368,
     mul_34_17_n_10369, mul_34_17_n_10370, mul_34_17_n_10371, mul_34_17_n_10372,
     mul_34_17_n_10373, mul_34_17_n_10374, mul_34_17_n_10375, mul_34_17_n_10376,
     mul_34_17_n_10377, mul_34_17_n_10378, mul_34_17_n_10379, mul_34_17_n_10380,
     mul_34_17_n_10381, mul_34_17_n_10382, mul_34_17_n_10383, mul_34_17_n_10384,
     mul_34_17_n_10385, mul_34_17_n_10386, mul_34_17_n_10387, mul_34_17_n_10388,
     mul_34_17_n_10389, mul_34_17_n_10390, mul_34_17_n_10391, mul_34_17_n_10392,
     mul_34_17_n_10393, mul_34_17_n_10394, mul_34_17_n_10395, mul_34_17_n_10396,
     mul_34_17_n_10397, mul_34_17_n_10398, mul_34_17_n_10399, mul_34_17_n_10400,
     mul_34_17_n_10401, mul_34_17_n_10402, mul_34_17_n_10403, mul_34_17_n_10404,
     mul_34_17_n_10405, mul_34_17_n_10406, mul_34_17_n_10407, mul_34_17_n_10408,
     mul_34_17_n_10409, mul_34_17_n_10410, mul_34_17_n_10411, mul_34_17_n_10412,
     mul_34_17_n_10413, mul_34_17_n_10414, mul_34_17_n_10415, mul_34_17_n_10416,
     mul_34_17_n_10417, mul_34_17_n_10418, mul_34_17_n_10419, mul_34_17_n_10420,
     mul_34_17_n_10421, mul_34_17_n_10422, mul_34_17_n_10423, mul_34_17_n_10424,
     mul_34_17_n_10425, mul_34_17_n_10426, mul_34_17_n_10427, mul_34_17_n_10428,
     mul_34_17_n_10429, mul_34_17_n_10430, mul_34_17_n_10431, mul_34_17_n_10432,
     mul_34_17_n_10433, mul_34_17_n_10434, mul_34_17_n_10435, mul_34_17_n_10436,
     mul_34_17_n_10437, mul_34_17_n_10438, mul_34_17_n_10439, mul_34_17_n_10440,
     mul_34_17_n_10441, mul_34_17_n_10442, mul_34_17_n_10443, mul_34_17_n_10444,
     mul_34_17_n_10445, mul_34_17_n_10446, mul_34_17_n_10447, mul_34_17_n_10448,
     mul_34_17_n_10449, mul_34_17_n_10450, mul_34_17_n_10451, mul_34_17_n_10452,
     mul_34_17_n_10453, mul_34_17_n_10454, mul_34_17_n_10455, mul_34_17_n_10456,
     mul_34_17_n_10457, mul_34_17_n_10458, mul_34_17_n_10459, mul_34_17_n_10460,
     mul_34_17_n_10461, mul_34_17_n_10462, mul_34_17_n_10463, mul_34_17_n_10464,
     mul_34_17_n_10465, mul_34_17_n_10466, mul_34_17_n_10467, mul_34_17_n_10468,
     mul_34_17_n_10469, mul_34_17_n_10470, mul_34_17_n_10471, mul_34_17_n_10472,
     mul_34_17_n_10473, mul_34_17_n_10474, mul_34_17_n_10475, mul_34_17_n_10476,
     mul_34_17_n_10477, mul_34_17_n_10478, mul_34_17_n_10479, mul_34_17_n_10480,
     mul_34_17_n_10481, mul_34_17_n_10482, mul_34_17_n_10483, mul_34_17_n_10484,
     mul_34_17_n_10485, mul_34_17_n_10486, mul_34_17_n_10487, mul_34_17_n_10488,
     mul_34_17_n_10489, mul_34_17_n_10490, mul_34_17_n_10491, mul_34_17_n_10492,
     mul_34_17_n_10493, mul_34_17_n_10494, mul_34_17_n_10495, mul_34_17_n_10496,
     mul_34_17_n_10497, mul_34_17_n_10498, mul_34_17_n_10499, mul_34_17_n_10500,
     mul_34_17_n_10501, mul_34_17_n_10502, mul_34_17_n_10503, mul_34_17_n_10504,
     mul_34_17_n_10505, mul_34_17_n_10506, mul_34_17_n_10507, mul_34_17_n_10508,
     mul_34_17_n_10509, mul_34_17_n_10510, mul_34_17_n_10511, mul_34_17_n_10512,
     mul_34_17_n_10513, mul_34_17_n_10514, mul_34_17_n_10515, mul_34_17_n_10516,
     mul_34_17_n_10517, mul_34_17_n_10518, mul_34_17_n_10519, mul_34_17_n_10520,
     mul_34_17_n_10521, mul_34_17_n_10522, mul_34_17_n_10523, mul_34_17_n_10524,
     mul_34_17_n_10525, mul_34_17_n_10526, mul_34_17_n_10527, mul_34_17_n_10528,
     mul_34_17_n_10529, mul_34_17_n_10530, mul_34_17_n_10531, mul_34_17_n_10532,
     mul_34_17_n_10533, mul_34_17_n_10534, mul_34_17_n_10535, mul_34_17_n_10536,
     mul_34_17_n_10537, mul_34_17_n_10538, mul_34_17_n_10539, mul_34_17_n_10540,
     mul_34_17_n_10541, mul_34_17_n_10542, mul_34_17_n_10543, mul_34_17_n_10544,
     mul_34_17_n_10545, mul_34_17_n_10546, mul_34_17_n_10547, mul_34_17_n_10548,
     mul_34_17_n_10549, mul_34_17_n_10550, mul_34_17_n_10551, mul_34_17_n_10552,
     mul_34_17_n_10553, mul_34_17_n_10554, mul_34_17_n_10555, mul_34_17_n_10556,
     mul_34_17_n_10557, mul_34_17_n_10558, mul_34_17_n_10559, mul_34_17_n_10560,
     mul_34_17_n_10561, mul_34_17_n_10562, mul_34_17_n_10563, mul_34_17_n_10564,
     mul_34_17_n_10565, mul_34_17_n_10566, mul_34_17_n_10567, mul_34_17_n_10568,
     mul_34_17_n_10569, mul_34_17_n_10570, mul_34_17_n_10571, mul_34_17_n_10572,
     mul_34_17_n_10573, mul_34_17_n_10574, mul_34_17_n_10575, mul_34_17_n_10576,
     mul_34_17_n_10577, mul_34_17_n_10578, mul_34_17_n_10579, mul_34_17_n_10580,
     mul_34_17_n_10581, mul_34_17_n_10582, mul_34_17_n_10583, mul_34_17_n_10584,
     mul_34_17_n_10585, mul_34_17_n_10586, mul_34_17_n_10587, mul_34_17_n_10588,
     mul_34_17_n_10589, mul_34_17_n_10590, mul_34_17_n_10591, mul_34_17_n_10592,
     mul_34_17_n_10593, mul_34_17_n_10594, mul_34_17_n_10595, mul_34_17_n_10596,
     mul_34_17_n_10597, mul_34_17_n_10598, mul_34_17_n_10599, mul_34_17_n_10600,
     mul_34_17_n_10601, mul_34_17_n_10602, mul_34_17_n_10603, mul_34_17_n_10604,
     mul_34_17_n_10605, mul_34_17_n_10606, mul_34_17_n_10607, mul_34_17_n_10608,
     mul_34_17_n_10609, mul_34_17_n_10610, mul_34_17_n_10611, mul_34_17_n_10612,
     mul_34_17_n_10613, mul_34_17_n_10614, mul_34_17_n_10615, mul_34_17_n_10616,
     mul_34_17_n_10617, mul_34_17_n_10618, mul_34_17_n_10619, mul_34_17_n_10620,
     mul_34_17_n_10621, mul_34_17_n_10622, mul_34_17_n_10623, mul_34_17_n_10624,
     mul_34_17_n_10625, mul_34_17_n_10626, mul_34_17_n_10627, mul_34_17_n_10628,
     mul_34_17_n_10629, mul_34_17_n_10630, mul_34_17_n_10631, mul_34_17_n_10632,
     mul_34_17_n_10633, mul_34_17_n_10634, mul_34_17_n_10635, mul_34_17_n_10636,
     mul_34_17_n_10637, mul_34_17_n_10638, mul_34_17_n_10639, mul_34_17_n_10640,
     mul_34_17_n_10641, mul_34_17_n_10642, mul_34_17_n_10643, mul_34_17_n_10644,
     mul_34_17_n_10645, mul_34_17_n_10646, mul_34_17_n_10647, mul_34_17_n_10648,
     mul_34_17_n_10649, mul_34_17_n_10650, mul_34_17_n_10651, mul_34_17_n_10652,
     mul_34_17_n_10653, mul_34_17_n_10654, mul_34_17_n_10655, mul_34_17_n_10656,
     mul_34_17_n_10657, mul_34_17_n_10658, mul_34_17_n_10659, mul_34_17_n_10660,
     mul_34_17_n_10661, mul_34_17_n_10662, mul_34_17_n_10663, mul_34_17_n_10664,
     mul_34_17_n_10665, mul_34_17_n_10666, mul_34_17_n_10667, mul_34_17_n_10668,
     mul_34_17_n_10669, mul_34_17_n_10670, mul_34_17_n_10671, mul_34_17_n_10672,
     mul_34_17_n_10673, mul_34_17_n_10674, mul_34_17_n_10675, mul_34_17_n_10676,
     mul_34_17_n_10677, mul_34_17_n_10678, mul_34_17_n_10679, mul_34_17_n_10680,
     mul_34_17_n_10681, mul_34_17_n_10682, mul_34_17_n_10683, mul_34_17_n_10684,
     mul_34_17_n_10685, mul_34_17_n_10686, mul_34_17_n_10687, mul_34_17_n_10688,
     mul_34_17_n_10689, mul_34_17_n_10690, mul_34_17_n_10691, mul_34_17_n_10692,
     mul_34_17_n_10693, mul_34_17_n_10694, mul_34_17_n_10695, mul_34_17_n_10696,
     mul_34_17_n_10697, mul_34_17_n_10698, mul_34_17_n_10699, mul_34_17_n_10700,
     mul_34_17_n_10701, mul_34_17_n_10702, mul_34_17_n_10703, mul_34_17_n_10704,
     mul_34_17_n_10705, mul_34_17_n_10706, mul_34_17_n_10707, mul_34_17_n_10708,
     mul_34_17_n_10709, mul_34_17_n_10710, mul_34_17_n_10711, mul_34_17_n_10712,
     mul_34_17_n_10713, mul_34_17_n_10714, mul_34_17_n_10715, mul_34_17_n_10716,
     mul_34_17_n_10717, mul_34_17_n_10718, mul_34_17_n_10719, mul_34_17_n_10720,
     mul_34_17_n_10721, mul_34_17_n_10722, mul_34_17_n_10723, mul_34_17_n_10724,
     mul_34_17_n_10725, mul_34_17_n_10726, mul_34_17_n_10727, mul_34_17_n_10728,
     mul_34_17_n_10729, mul_34_17_n_10730, mul_34_17_n_10731, mul_34_17_n_10732,
     mul_34_17_n_10733, mul_34_17_n_10734, mul_34_17_n_10735, mul_34_17_n_10736,
     mul_34_17_n_10737, mul_34_17_n_10738, mul_34_17_n_10739, mul_34_17_n_10740,
     mul_34_17_n_10741, mul_34_17_n_10742, mul_34_17_n_10743, mul_34_17_n_10744,
     mul_34_17_n_10745, mul_34_17_n_10746, mul_34_17_n_10747, mul_34_17_n_10748,
     mul_34_17_n_10749, mul_34_17_n_10750, mul_34_17_n_10751, mul_34_17_n_10752,
     mul_34_17_n_10753, mul_34_17_n_10754, mul_34_17_n_10755, mul_34_17_n_10756,
     mul_34_17_n_10757, mul_34_17_n_10758, mul_34_17_n_10759, mul_34_17_n_10760,
     mul_34_17_n_10761, mul_34_17_n_10762, mul_34_17_n_10763, mul_34_17_n_10764,
     mul_34_17_n_10765, mul_34_17_n_10766, mul_34_17_n_10767, mul_34_17_n_10768,
     mul_34_17_n_10769, mul_34_17_n_10770, mul_34_17_n_10771, mul_34_17_n_10772,
     mul_34_17_n_10773, mul_34_17_n_10774, mul_34_17_n_10775, mul_34_17_n_10776,
     mul_34_17_n_10777, mul_34_17_n_10778, mul_34_17_n_10779, mul_34_17_n_10780,
     mul_34_17_n_10781, mul_34_17_n_10782, mul_34_17_n_10783, mul_34_17_n_10784,
     mul_34_17_n_10785, mul_34_17_n_10786, mul_34_17_n_10787, mul_34_17_n_10788,
     mul_34_17_n_10789, mul_34_17_n_10790, mul_34_17_n_10791, mul_34_17_n_10792,
     mul_34_17_n_10793, mul_34_17_n_10794, mul_34_17_n_10795, mul_34_17_n_10796,
     mul_34_17_n_10797, mul_34_17_n_10798, mul_34_17_n_10799, mul_34_17_n_10800,
     mul_34_17_n_10801, mul_34_17_n_10802, mul_34_17_n_10803, mul_34_17_n_10804,
     mul_34_17_n_10805, mul_34_17_n_10806, mul_34_17_n_10807, mul_34_17_n_10808,
     mul_34_17_n_10809, mul_34_17_n_10810, mul_34_17_n_10811, mul_34_17_n_10812,
     mul_34_17_n_10813, mul_34_17_n_10814, mul_34_17_n_10815, mul_34_17_n_10816,
     mul_34_17_n_10817, mul_34_17_n_10818, mul_34_17_n_10819, mul_34_17_n_10820,
     mul_34_17_n_10821, mul_34_17_n_10822, mul_34_17_n_10823, mul_34_17_n_10824,
     mul_34_17_n_10825, mul_34_17_n_10826, mul_34_17_n_10827, mul_34_17_n_10828,
     mul_34_17_n_10829, mul_34_17_n_10830, mul_34_17_n_10831, mul_34_17_n_10832,
     mul_34_17_n_10833, mul_34_17_n_10834, mul_34_17_n_10835, mul_34_17_n_10836,
     mul_34_17_n_10837, mul_34_17_n_10838, mul_34_17_n_10839, mul_34_17_n_10840,
     mul_34_17_n_10841, mul_34_17_n_10842, mul_34_17_n_10843, mul_34_17_n_10844,
     mul_34_17_n_10845, mul_34_17_n_10846, mul_34_17_n_10847, mul_34_17_n_10848,
     mul_34_17_n_10849, mul_34_17_n_10850, mul_34_17_n_10851, mul_34_17_n_10852,
     mul_34_17_n_10853, mul_34_17_n_10854, mul_34_17_n_10855, mul_34_17_n_10856,
     mul_34_17_n_10857, mul_34_17_n_10858, mul_34_17_n_10859, mul_34_17_n_10860,
     mul_34_17_n_10861, mul_34_17_n_10862, mul_34_17_n_10863, mul_34_17_n_10864,
     mul_34_17_n_10865, mul_34_17_n_10866, mul_34_17_n_10867, mul_34_17_n_10868,
     mul_34_17_n_10869, mul_34_17_n_10870, mul_34_17_n_10871, mul_34_17_n_10872,
     mul_34_17_n_10873, mul_34_17_n_10874, mul_34_17_n_10875, mul_34_17_n_10876,
     mul_34_17_n_10877, mul_34_17_n_10878, mul_34_17_n_10879, mul_34_17_n_10880,
     mul_34_17_n_10881, mul_34_17_n_10882, mul_34_17_n_10883, mul_34_17_n_10884,
     mul_34_17_n_10885, mul_34_17_n_10886, mul_34_17_n_10887, mul_34_17_n_10888,
     mul_34_17_n_10889, mul_34_17_n_10890, mul_34_17_n_10891, mul_34_17_n_10892,
     mul_34_17_n_10893, mul_34_17_n_10894, mul_34_17_n_10895, mul_34_17_n_10896,
     mul_34_17_n_10897, mul_34_17_n_10898, mul_34_17_n_10899, mul_34_17_n_10900,
     mul_34_17_n_10901, mul_34_17_n_10902, mul_34_17_n_10903, mul_34_17_n_10904,
     mul_34_17_n_10905, mul_34_17_n_10906, mul_34_17_n_10907, mul_34_17_n_10908,
     mul_34_17_n_10909, mul_34_17_n_10910, mul_34_17_n_10911, mul_34_17_n_10912,
     mul_34_17_n_10913, mul_34_17_n_10914, mul_34_17_n_10915, mul_34_17_n_10916,
     mul_34_17_n_10917, mul_34_17_n_10918, mul_34_17_n_10919, mul_34_17_n_10920,
     mul_34_17_n_10921, mul_34_17_n_10922, mul_34_17_n_10923, mul_34_17_n_10924,
     mul_34_17_n_10925, mul_34_17_n_10926, mul_34_17_n_10927, mul_34_17_n_10928,
     mul_34_17_n_10929, mul_34_17_n_10930, mul_34_17_n_10931, mul_34_17_n_10932,
     mul_34_17_n_10933, mul_34_17_n_10934, mul_34_17_n_10935, mul_34_17_n_10936,
     mul_34_17_n_10937, mul_34_17_n_10938, mul_34_17_n_10939, mul_34_17_n_10940,
     mul_34_17_n_10941, mul_34_17_n_10942, mul_34_17_n_10943, mul_34_17_n_10944,
     mul_34_17_n_10945, mul_34_17_n_10946, mul_34_17_n_10947, mul_34_17_n_10948,
     mul_34_17_n_10949, mul_34_17_n_10950, mul_34_17_n_10951, mul_34_17_n_10952,
     mul_34_17_n_10953, mul_34_17_n_10954, mul_34_17_n_10955, mul_34_17_n_10956,
     mul_34_17_n_10957, mul_34_17_n_10958, mul_34_17_n_10959, mul_34_17_n_10960,
     mul_34_17_n_10961, mul_34_17_n_10962, mul_34_17_n_10963, mul_34_17_n_10964,
     mul_34_17_n_10965, mul_34_17_n_10966, mul_34_17_n_10967, mul_34_17_n_10968,
     mul_34_17_n_10969, mul_34_17_n_10970, mul_34_17_n_10971, mul_34_17_n_10972,
     mul_34_17_n_10973, mul_34_17_n_10974, mul_34_17_n_10975, mul_34_17_n_10976,
     mul_34_17_n_10977, mul_34_17_n_10978, mul_34_17_n_10979, mul_34_17_n_10980,
     mul_34_17_n_10981, mul_34_17_n_10982, mul_34_17_n_10983, mul_34_17_n_10984,
     mul_34_17_n_10985, mul_34_17_n_10986, mul_34_17_n_10987, mul_34_17_n_10988,
     mul_34_17_n_10989, mul_34_17_n_10990, mul_34_17_n_10991, mul_34_17_n_10992,
     mul_34_17_n_10993, mul_34_17_n_10994, mul_34_17_n_10995, mul_34_17_n_10996,
     mul_34_17_n_10997, mul_34_17_n_10998, mul_34_17_n_10999, mul_34_17_n_11000,
     mul_34_17_n_11001, mul_34_17_n_11002, mul_34_17_n_11003, mul_34_17_n_11004,
     mul_34_17_n_11005, mul_34_17_n_11006, mul_34_17_n_11007, mul_34_17_n_11008,
     mul_34_17_n_11009, mul_34_17_n_11010, mul_34_17_n_11011, mul_34_17_n_11012,
     mul_34_17_n_11013, mul_34_17_n_11014, mul_34_17_n_11015, mul_34_17_n_11016,
     mul_34_17_n_11017, mul_34_17_n_11018, mul_34_17_n_11019, mul_34_17_n_11020,
     mul_34_17_n_11021, mul_34_17_n_11022, mul_34_17_n_11023, mul_34_17_n_11024,
     mul_34_17_n_11025, mul_34_17_n_11026, mul_34_17_n_11027, mul_34_17_n_11028,
     mul_34_17_n_11029, mul_34_17_n_11030, mul_34_17_n_11031, mul_34_17_n_11032,
     mul_34_17_n_11033, mul_34_17_n_11034, mul_34_17_n_11035, mul_34_17_n_11036,
     mul_34_17_n_11037, mul_34_17_n_11038, mul_34_17_n_11039, mul_34_17_n_11040,
     mul_34_17_n_11041, mul_34_17_n_11042, mul_34_17_n_11043, mul_34_17_n_11044,
     mul_34_17_n_11045, mul_34_17_n_11046, mul_34_17_n_11047, mul_34_17_n_11048,
     mul_34_17_n_11049, mul_34_17_n_11050, mul_34_17_n_11247, mul_34_17_n_11248,
     mul_34_17_n_11251, mul_34_17_n_11252, mul_34_17_n_11253, mul_34_17_n_11272,
     mul_34_17_n_11273, mul_34_17_n_11274, mul_34_17_n_11275, mul_34_17_n_11276,
     mul_34_17_n_11277, mul_34_17_n_11278, mul_34_17_n_11279, mul_34_17_n_11280,
     mul_34_17_n_11281, mul_34_17_n_11282, mul_34_17_n_11283, mul_34_17_n_11284,
     mul_34_17_n_11285, mul_34_17_n_11286, mul_34_17_n_11287, mul_34_17_n_11288,
     mul_34_17_n_11289, mul_34_17_n_11290, mul_34_17_n_11291, mul_34_17_n_11292,
     mul_34_17_n_11293, mul_34_17_n_11294, mul_34_17_n_11295, mul_34_17_n_11296,
     mul_34_17_n_11297, mul_34_17_n_11298, mul_34_17_n_11299, mul_34_17_n_11300,
     mul_34_17_n_11301, mul_34_17_n_11302, mul_34_17_n_11303, mul_34_17_n_11304,
     mul_34_17_n_11305, mul_34_17_n_11306, mul_34_17_n_11307, mul_34_17_n_11308,
     mul_34_17_n_11309, mul_34_17_n_11310, mul_34_17_n_11311, mul_34_17_n_11312,
     mul_34_17_n_11313, mul_34_17_n_11314, mul_34_17_n_11315, mul_34_17_n_11316,
     mul_34_17_n_11317, mul_34_17_n_11318, mul_34_17_n_11319, mul_34_17_n_11320,
     mul_34_17_n_11321, mul_34_17_n_11322, mul_34_17_n_11323, mul_34_17_n_11324,
     mul_34_17_n_11325, mul_34_17_n_11326, mul_34_17_n_11327, mul_34_17_n_11328,
     mul_34_17_n_11329, mul_34_17_n_11330, mul_34_17_n_11331, mul_34_17_n_11332,
     mul_34_17_n_11333, mul_34_17_n_11334, mul_34_17_n_11335, mul_34_17_n_11336,
     mul_34_17_n_11337, mul_34_17_n_11338, mul_34_17_n_11339, mul_34_17_n_11340,
     mul_34_17_n_11341, mul_34_17_n_11342, mul_34_17_n_11343, mul_34_17_n_11344,
     mul_34_17_n_11345, mul_34_17_n_11346, mul_34_17_n_11347, mul_34_17_n_11348,
     mul_34_17_n_11349, mul_34_17_n_11350, mul_34_17_n_11351, mul_34_17_n_11352,
     mul_34_17_n_11353, mul_34_17_n_11354, mul_34_17_n_11355, mul_34_17_n_11356,
     mul_34_17_n_11357, mul_34_17_n_11358, mul_34_17_n_11359, mul_34_17_n_11360,
     mul_34_17_n_11361, mul_34_17_n_11362, mul_34_17_n_11363, mul_34_17_n_11364,
     mul_34_17_n_11365, mul_34_17_n_11366, mul_34_17_n_11367, mul_34_17_n_11368,
     mul_34_17_n_11369, mul_34_17_n_11370, mul_34_17_n_11371, mul_34_17_n_11372,
     mul_34_17_n_11373, mul_34_17_n_11374, mul_34_17_n_11375, mul_34_17_n_11376,
     mul_34_17_n_11377, mul_34_17_n_11378, mul_34_17_n_11379, mul_34_17_n_11380,
     mul_34_17_n_11381, mul_34_17_n_11382, mul_34_17_n_11383, mul_34_17_n_11384,
     mul_34_17_n_11385, mul_34_17_n_11386, mul_34_17_n_11387, mul_34_17_n_11388,
     mul_34_17_n_11389, mul_34_17_n_11390, mul_34_17_n_11391, mul_34_17_n_11392,
     mul_34_17_n_11393, mul_34_17_n_11394, mul_34_17_n_11395, mul_34_17_n_11396,
     mul_34_17_n_11397, mul_34_17_n_11398, mul_34_17_n_11399, mul_34_17_n_11400,
     mul_34_17_n_11401, mul_34_17_n_11402, mul_34_17_n_11403, mul_34_17_n_11404,
     mul_34_17_n_11405, mul_34_17_n_11406, mul_34_17_n_11407, mul_34_17_n_11408,
     mul_34_17_n_11409, mul_34_17_n_11410, mul_34_17_n_11411, mul_34_17_n_11412,
     mul_34_17_n_11413, mul_34_17_n_11414, mul_34_17_n_11415, mul_34_17_n_11416,
     mul_34_17_n_11417, mul_34_17_n_11418, mul_34_17_n_11419, mul_34_17_n_11420,
     mul_34_17_n_11421, mul_34_17_n_11422, mul_34_17_n_11423, mul_34_17_n_11424,
     mul_34_17_n_11425, mul_34_17_n_11426, mul_34_17_n_11427, mul_34_17_n_11428,
     mul_34_17_n_11429, mul_34_17_n_11430, mul_34_17_n_11431, mul_34_17_n_11432,
     mul_34_17_n_11433, mul_34_17_n_11434, mul_34_17_n_11435, mul_34_17_n_11436,
     mul_34_17_n_11437, mul_34_17_n_11438, mul_34_17_n_11439, mul_34_17_n_11440,
     mul_34_17_n_11441, mul_34_17_n_11442, mul_34_17_n_11443, mul_34_17_n_11444,
     mul_34_17_n_11445, mul_34_17_n_11446, mul_34_17_n_11447, mul_34_17_n_11448,
     mul_34_17_n_11449, mul_34_17_n_11450, mul_34_17_n_11451, mul_34_17_n_11452,
     mul_34_17_n_11453, mul_34_17_n_11454, mul_34_17_n_11455, mul_34_17_n_11456,
     mul_34_17_n_11457, mul_34_17_n_11458, mul_34_17_n_11459, mul_34_17_n_11460,
     mul_34_17_n_11461, mul_34_17_n_11462, mul_34_17_n_11463, mul_34_17_n_11464,
     mul_34_17_n_11465, mul_34_17_n_11466, mul_34_17_n_11467, mul_34_17_n_11468,
     mul_34_17_n_11469, mul_34_17_n_11470, mul_34_17_n_11471, mul_34_17_n_11472,
     mul_34_17_n_11473, mul_34_17_n_11474, mul_34_17_n_11475, mul_34_17_n_11476,
     mul_34_17_n_11477, mul_34_17_n_11478, mul_34_17_n_11479, mul_34_17_n_11480,
     mul_34_17_n_11481, mul_34_17_n_11482, mul_34_17_n_11483, mul_34_17_n_11484,
     mul_34_17_n_11485, mul_34_17_n_11486, mul_34_17_n_11487, mul_34_17_n_11488,
     mul_34_17_n_11489, mul_34_17_n_11490, mul_34_17_n_11491, mul_34_17_n_11492,
     mul_34_17_n_11493, mul_34_17_n_11494, mul_34_17_n_11495, mul_34_17_n_11496,
     mul_34_17_n_11497, mul_34_17_n_11498, mul_34_17_n_11499, mul_34_17_n_11500,
     mul_34_17_n_11501, mul_34_17_n_11502, mul_34_17_n_11503, mul_34_17_n_11504,
     mul_34_17_n_11513, mul_34_17_n_11514, mul_34_17_n_11515, mul_34_17_n_11516,
     mul_34_17_n_11517, mul_34_17_n_11518, mul_34_17_n_11519, mul_34_17_n_11520,
     mul_34_17_n_11521, mul_34_17_n_11522, mul_34_17_n_11523, mul_34_17_n_11524,
     mul_34_17_n_11525, mul_34_17_n_11526, mul_34_17_n_11527, mul_34_17_n_11528,
     mul_34_17_n_11529, mul_34_17_n_11530, mul_34_17_n_11531, mul_34_17_n_11532,
     mul_34_17_n_11533, mul_34_17_n_11534, mul_34_17_n_11535, mul_34_17_n_11536,
     mul_34_17_n_11537, mul_34_17_n_11538, mul_34_17_n_11539, mul_34_17_n_11540,
     mul_34_17_n_11541, mul_34_17_n_11542, mul_34_17_n_11543, mul_34_17_n_11544,
     mul_34_17_n_11545, mul_34_17_n_11546, mul_34_17_n_11547, mul_34_17_n_11548,
     mul_34_17_n_11549, mul_34_17_n_11550, mul_34_17_n_11551, mul_34_17_n_11552,
     mul_34_17_n_11553, mul_34_17_n_11554, mul_34_17_n_11555, mul_34_17_n_11556,
     mul_34_17_n_11557, mul_34_17_n_11558, mul_34_17_n_11559, mul_34_17_n_11560,
     mul_34_17_n_11561, mul_34_17_n_11562, mul_34_17_n_11563, mul_34_17_n_11564,
     mul_34_17_n_11565, mul_34_17_n_11566, mul_34_17_n_11567, mul_34_17_n_11568,
     mul_34_17_n_11569, mul_34_17_n_11570, mul_34_17_n_11571, mul_34_17_n_11572,
     mul_34_17_n_11573, mul_34_17_n_11574, mul_34_17_n_11575, mul_34_17_n_11576,
     mul_34_17_n_11577, mul_34_17_n_11578, mul_34_17_n_11579, mul_34_17_n_11580,
     mul_34_17_n_11581, mul_34_17_n_11582, mul_34_17_n_11583, mul_34_17_n_11584,
     mul_34_17_n_11585, mul_34_17_n_11586, mul_34_17_n_11587, mul_34_17_n_11588,
     mul_34_17_n_11589, mul_34_17_n_11590, mul_34_17_n_11591, mul_34_17_n_11592,
     mul_34_17_n_11593, mul_34_17_n_11595, mul_34_17_n_11596, mul_34_17_n_11597,
     mul_34_17_n_11598, mul_34_17_n_11599, mul_34_17_n_11600, mul_34_17_n_11601,
     mul_34_17_n_11602, mul_34_17_n_11603, mul_34_17_n_11604, mul_34_17_n_11605,
     mul_34_17_n_11606, mul_34_17_n_11607, mul_34_17_n_11608, mul_34_17_n_11609,
     mul_34_17_n_11610, mul_34_17_n_11611, mul_34_17_n_11612, mul_34_17_n_11613,
     mul_34_17_n_11614, mul_34_17_n_11615, mul_34_17_n_11616, mul_34_17_n_11617,
     mul_34_17_n_11618, mul_34_17_n_11619, mul_34_17_n_11620, mul_34_17_n_11621,
     mul_34_17_n_11622, mul_34_17_n_11623, mul_34_17_n_11624, mul_34_17_n_11625,
     mul_34_17_n_11626, mul_34_17_n_11627, mul_34_17_n_11628, mul_34_17_n_11629,
     mul_34_17_n_11630, mul_34_17_n_11631, mul_34_17_n_11632, mul_34_17_n_11633,
     mul_34_17_n_11634, mul_34_17_n_11635, mul_34_17_n_11636, mul_34_17_n_11637,
     mul_34_17_n_11638, mul_34_17_n_11639, mul_34_17_n_11640, mul_34_17_n_11641,
     mul_34_17_n_11642, mul_34_17_n_11643, mul_34_17_n_11644, mul_34_17_n_11645,
     mul_34_17_n_11646, mul_34_17_n_11648, mul_34_17_n_11649, mul_34_17_n_11651,
     mul_34_17_n_11652, mul_34_17_n_11653, mul_34_17_n_11658, mul_34_17_n_11659,
     mul_34_17_n_11660, mul_34_17_n_11662, mul_34_17_n_11663, mul_34_17_n_11665,
     mul_34_17_n_11666, mul_34_17_n_11672, mul_34_17_n_11673, mul_34_17_n_11675,
     mul_34_17_n_11676, mul_34_17_n_11678, mul_34_17_n_11679, mul_34_17_n_11680,
     mul_34_17_n_11682, mul_34_17_n_11683, mul_34_17_n_11685, mul_34_17_n_11686,
     mul_34_17_n_11693, mul_34_17_n_11694, mul_34_17_n_11696, mul_34_17_n_11697,
     asc001_0_, asc001_1_, asc001_2_, asc001_3_, asc001_4_, asc001_5_, asc001_6_,
     asc001_7_, asc001_8_, asc001_9_, asc001_10_, asc001_11_, asc001_12_,
     asc001_13_, asc001_14_, asc001_15_, asc001_16_, asc001_17_, asc001_18_,
     asc001_19_, asc001_20_, asc001_21_, asc001_22_, asc001_23_, asc001_24_,
     asc001_25_, asc001_26_, asc001_27_, asc001_28_, asc001_29_, asc001_30_,
     asc001_31_, asc001_32_, asc001_33_, asc001_34_, asc001_35_, asc001_36_,
     asc001_37_, asc001_38_, asc001_39_, asc001_40_, asc001_41_, asc001_42_,
     asc001_43_, asc001_44_, asc001_45_, asc001_46_, asc001_47_, asc001_48_,
     asc001_49_, asc001_50_, asc001_51_, asc001_52_, asc001_53_, asc001_54_,
     asc001_55_, asc001_56_, asc001_57_, asc001_58_, asc001_59_, asc001_60_,
     asc001_61_, asc001_62_, asc001_63_, asc001_64_, asc001_65_, asc001_66_,
     asc001_67_, asc001_68_, asc001_69_, asc001_70_, asc001_71_, asc001_72_,
     asc001_73_, asc001_74_, asc001_75_, asc001_76_, asc001_77_, asc001_78_,
     asc001_79_, asc001_80_, asc001_81_, asc001_82_, asc001_83_, asc001_84_,
     asc001_85_, in;
assign {out1[85]} = asc001_85_;
assign {out1[84]} = asc001_84_;
assign {out1[83]} = asc001_83_;
assign {out1[82]} = asc001_82_;
assign {out1[81]} = asc001_81_;
assign {out1[80]} = asc001_80_;
assign {out1[79]} = asc001_79_;
assign {out1[78]} = asc001_78_;
assign {out1[77]} = asc001_77_;
assign {out1[76]} = asc001_76_;
assign {out1[75]} = asc001_75_;
assign {out1[74]} = asc001_74_;
assign {out1[73]} = asc001_73_;
assign {out1[72]} = asc001_72_;
assign {out1[71]} = asc001_71_;
assign {out1[70]} = asc001_70_;
assign {out1[69]} = asc001_69_;
assign {out1[68]} = asc001_68_;
assign {out1[67]} = asc001_67_;
assign {out1[66]} = asc001_66_;
assign {out1[65]} = asc001_65_;
assign {out1[64]} = asc001_64_;
assign {out1[63]} = asc001_63_;
assign {out1[62]} = asc001_62_;
assign {out1[61]} = asc001_61_;
assign {out1[60]} = asc001_60_;
assign {out1[59]} = asc001_59_;
assign {out1[58]} = asc001_58_;
assign {out1[57]} = asc001_57_;
assign {out1[56]} = asc001_56_;
assign {out1[55]} = asc001_55_;
assign {out1[54]} = asc001_54_;
assign {out1[53]} = asc001_53_;
assign {out1[52]} = asc001_52_;
assign {out1[51]} = asc001_51_;
assign {out1[50]} = asc001_50_;
assign {out1[49]} = asc001_49_;
assign {out1[48]} = asc001_48_;
assign {out1[47]} = asc001_47_;
assign {out1[46]} = asc001_46_;
assign {out1[45]} = asc001_45_;
assign {out1[44]} = asc001_44_;
assign {out1[43]} = asc001_43_;
assign {out1[42]} = asc001_42_;
assign {out1[41]} = asc001_41_;
assign {out1[40]} = asc001_40_;
assign {out1[39]} = asc001_39_;
assign {out1[38]} = asc001_38_;
assign {out1[37]} = asc001_37_;
assign {out1[36]} = asc001_36_;
assign {out1[35]} = asc001_35_;
assign {out1[34]} = asc001_34_;
assign {out1[33]} = asc001_33_;
assign {out1[32]} = asc001_32_;
assign {out1[31]} = asc001_31_;
assign {out1[30]} = asc001_30_;
assign {out1[29]} = asc001_29_;
assign {out1[28]} = asc001_28_;
assign {out1[27]} = asc001_27_;
assign {out1[26]} = asc001_26_;
assign {out1[25]} = asc001_25_;
assign {out1[24]} = asc001_24_;
assign {out1[23]} = asc001_23_;
assign {out1[22]} = asc001_22_;
assign {out1[21]} = asc001_21_;
assign {out1[20]} = asc001_20_;
assign {out1[19]} = asc001_19_;
assign {out1[18]} = asc001_18_;
assign {out1[17]} = asc001_17_;
assign {out1[16]} = asc001_16_;
assign {out1[15]} = asc001_15_;
assign {out1[14]} = asc001_14_;
assign {out1[13]} = asc001_13_;
assign {out1[12]} = asc001_12_;
assign {out1[11]} = asc001_11_;
assign {out1[10]} = asc001_10_;
assign {out1[9]} = asc001_9_;
assign {out1[8]} = asc001_8_;
assign {out1[7]} = asc001_7_;
assign {out1[6]} = asc001_6_;
assign {out1[5]} = asc001_5_;
assign {out1[4]} = asc001_4_;
assign {out1[3]} = asc001_3_;
assign {out1[2]} = asc001_2_;
assign {out1[1]} = asc001_1_;
assign {out1[0]} = asc001_0_;
 reg mul_34_17_retime_s1_1_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_1_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_1_reg_reg_IQ <= mul_34_17_n_9729;
     end
 assign mul_34_17_n_10825 = mul_34_17_retime_s1_1_reg_reg_IQ;
 reg mul_34_17_retime_s1_2_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_2_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_2_reg_reg_IQ <= mul_34_17_n_10175;
     end
 assign mul_34_17_n_10826 = mul_34_17_retime_s1_2_reg_reg_IQ;
 reg mul_34_17_retime_s1_3_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_3_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_3_reg_reg_IQ <= mul_34_17_n_10269;
     end
 assign mul_34_17_n_10827 = mul_34_17_retime_s1_3_reg_reg_IQ;
 reg mul_34_17_retime_s1_4_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_4_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_4_reg_reg_IQ <= mul_34_17_n_10124;
     end
 assign mul_34_17_n_10828 = mul_34_17_retime_s1_4_reg_reg_IQ;
 reg mul_34_17_retime_s1_5_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_5_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_5_reg_reg_IQ <= mul_34_17_n_10072;
     end
 assign mul_34_17_n_10829 = mul_34_17_retime_s1_5_reg_reg_IQ;
 reg mul_34_17_retime_s1_6_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_6_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_6_reg_reg_IQ <= mul_34_17_n_10169;
     end
 assign mul_34_17_n_10830 = mul_34_17_retime_s1_6_reg_reg_IQ;
 reg mul_34_17_retime_s1_7_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_7_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_7_reg_reg_IQ <= mul_34_17_n_10280;
     end
 assign mul_34_17_n_10831 = mul_34_17_retime_s1_7_reg_reg_IQ;
 reg mul_34_17_retime_s1_8_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_8_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_8_reg_reg_IQ <= mul_34_17_n_10224;
     end
 assign mul_34_17_n_10832 = mul_34_17_retime_s1_8_reg_reg_IQ;
 reg mul_34_17_retime_s1_9_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_9_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_9_reg_reg_IQ <= mul_34_17_n_9403;
     end
 assign mul_34_17_n_10833 = mul_34_17_retime_s1_9_reg_reg_IQ;
 reg mul_34_17_retime_s1_10_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_10_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_10_reg_reg_IQ <= mul_34_17_n_9919;
     end
 assign mul_34_17_n_10834 = mul_34_17_retime_s1_10_reg_reg_IQ;
 reg mul_34_17_retime_s1_11_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_11_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_11_reg_reg_IQ <= mul_34_17_n_10207;
     end
 assign mul_34_17_n_10835 = mul_34_17_retime_s1_11_reg_reg_IQ;
 reg mul_34_17_retime_s1_12_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_12_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_12_reg_reg_IQ <= mul_34_17_n_9875;
     end
 assign mul_34_17_n_10836 = mul_34_17_retime_s1_12_reg_reg_IQ;
 reg mul_34_17_retime_s1_13_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_13_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_13_reg_reg_IQ <= mul_34_17_n_9877;
     end
 assign mul_34_17_n_10837 = mul_34_17_retime_s1_13_reg_reg_IQ;
 reg mul_34_17_retime_s1_14_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_14_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_14_reg_reg_IQ <= mul_34_17_n_323;
     end
 assign mul_34_17_n_10838 = mul_34_17_retime_s1_14_reg_reg_IQ;
 reg mul_34_17_retime_s1_15_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_15_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_15_reg_reg_IQ <= mul_34_17_n_10281;
     end
 assign mul_34_17_n_10839 = mul_34_17_retime_s1_15_reg_reg_IQ;
 reg mul_34_17_retime_s1_16_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_16_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_16_reg_reg_IQ <= mul_34_17_n_9913;
     end
 assign mul_34_17_n_10840 = mul_34_17_retime_s1_16_reg_reg_IQ;
 reg mul_34_17_retime_s1_17_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_17_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_17_reg_reg_IQ <= mul_34_17_n_10206;
     end
 assign mul_34_17_n_10841 = mul_34_17_retime_s1_17_reg_reg_IQ;
 reg mul_34_17_retime_s1_18_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_18_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_18_reg_reg_IQ <= mul_34_17_n_10238;
     end
 assign mul_34_17_n_11248 = mul_34_17_retime_s1_18_reg_reg_IQ;
 reg mul_34_17_retime_s1_19_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_19_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_19_reg_reg_IQ <= mul_34_17_n_10077;
     end
 assign mul_34_17_n_10842 = mul_34_17_retime_s1_19_reg_reg_IQ;
 reg mul_34_17_retime_s1_20_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_20_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_20_reg_reg_IQ <= mul_34_17_n_10240;
     end
 assign mul_34_17_n_10843 = mul_34_17_retime_s1_20_reg_reg_IQ;
 reg mul_34_17_retime_s1_21_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_21_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_21_reg_reg_IQ <= mul_34_17_n_292;
     end
 assign mul_34_17_n_10844 = mul_34_17_retime_s1_21_reg_reg_IQ;
 reg mul_34_17_retime_s1_22_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_22_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_22_reg_reg_IQ <= mul_34_17_n_10078;
     end
 assign mul_34_17_n_10845 = mul_34_17_retime_s1_22_reg_reg_IQ;
 reg mul_34_17_retime_s1_23_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_23_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_23_reg_reg_IQ <= mul_34_17_n_10041;
     end
 assign mul_34_17_n_10846 = mul_34_17_retime_s1_23_reg_reg_IQ;
 reg mul_34_17_retime_s1_24_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_24_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_24_reg_reg_IQ <= mul_34_17_n_10259;
     end
 assign mul_34_17_n_10847 = mul_34_17_retime_s1_24_reg_reg_IQ;
 reg mul_34_17_retime_s1_25_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_25_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_25_reg_reg_IQ <= mul_34_17_n_10141;
     end
 assign mul_34_17_n_10848 = mul_34_17_retime_s1_25_reg_reg_IQ;
 reg mul_34_17_retime_s1_26_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_26_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_26_reg_reg_IQ <= mul_34_17_n_10115;
     end
 assign mul_34_17_n_10849 = mul_34_17_retime_s1_26_reg_reg_IQ;
 reg mul_34_17_retime_s1_27_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_27_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_27_reg_reg_IQ <= mul_34_17_n_10128;
     end
 assign mul_34_17_n_10850 = mul_34_17_retime_s1_27_reg_reg_IQ;
 reg mul_34_17_retime_s1_28_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_28_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_28_reg_reg_IQ <= mul_34_17_n_8703;
     end
 assign mul_34_17_n_10851 = mul_34_17_retime_s1_28_reg_reg_IQ;
 reg mul_34_17_retime_s1_29_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_29_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_29_reg_reg_IQ <= mul_34_17_n_9515;
     end
 assign mul_34_17_n_10852 = mul_34_17_retime_s1_29_reg_reg_IQ;
 reg mul_34_17_retime_s1_30_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_30_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_30_reg_reg_IQ <= mul_34_17_n_10258;
     end
 assign mul_34_17_n_10853 = mul_34_17_retime_s1_30_reg_reg_IQ;
 reg mul_34_17_retime_s1_31_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_31_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_31_reg_reg_IQ <= mul_34_17_n_10230;
     end
 assign mul_34_17_n_11247 = mul_34_17_retime_s1_31_reg_reg_IQ;
 reg mul_34_17_retime_s1_32_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_32_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_32_reg_reg_IQ <= mul_34_17_n_342;
     end
 assign mul_34_17_n_10854 = mul_34_17_retime_s1_32_reg_reg_IQ;
 reg mul_34_17_retime_s1_33_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_33_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_33_reg_reg_IQ <= mul_34_17_n_315;
     end
 assign mul_34_17_n_10855 = mul_34_17_retime_s1_33_reg_reg_IQ;
 reg mul_34_17_retime_s1_34_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_34_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_34_reg_reg_IQ <= mul_34_17_n_10236;
     end
 assign mul_34_17_n_10856 = mul_34_17_retime_s1_34_reg_reg_IQ;
 reg mul_34_17_retime_s1_35_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_35_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_35_reg_reg_IQ <= mul_34_17_n_10278;
     end
 assign mul_34_17_n_10857 = mul_34_17_retime_s1_35_reg_reg_IQ;
 reg mul_34_17_retime_s1_36_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_36_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_36_reg_reg_IQ <= mul_34_17_n_10076;
     end
 assign mul_34_17_n_10858 = mul_34_17_retime_s1_36_reg_reg_IQ;
 reg mul_34_17_retime_s1_37_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_37_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_37_reg_reg_IQ <= mul_34_17_n_10205;
     end
 assign mul_34_17_n_10859 = mul_34_17_retime_s1_37_reg_reg_IQ;
 reg mul_34_17_retime_s1_38_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_38_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_38_reg_reg_IQ <= mul_34_17_n_10075;
     end
 assign mul_34_17_n_10860 = mul_34_17_retime_s1_38_reg_reg_IQ;
 reg mul_34_17_retime_s1_39_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_39_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_39_reg_reg_IQ <= mul_34_17_n_10034;
     end
 assign mul_34_17_n_10861 = mul_34_17_retime_s1_39_reg_reg_IQ;
 reg mul_34_17_retime_s1_40_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_40_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_40_reg_reg_IQ <= mul_34_17_n_10227;
     end
 assign mul_34_17_n_10862 = mul_34_17_retime_s1_40_reg_reg_IQ;
 reg mul_34_17_retime_s1_41_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_41_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_41_reg_reg_IQ <= mul_34_17_n_340;
     end
 assign mul_34_17_n_10863 = mul_34_17_retime_s1_41_reg_reg_IQ;
 reg mul_34_17_retime_s1_42_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_42_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_42_reg_reg_IQ <= mul_34_17_n_10132;
     end
 assign mul_34_17_n_10864 = mul_34_17_retime_s1_42_reg_reg_IQ;
 reg mul_34_17_retime_s1_43_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_43_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_43_reg_reg_IQ <= mul_34_17_n_9834;
     end
 assign mul_34_17_n_10865 = mul_34_17_retime_s1_43_reg_reg_IQ;
 reg mul_34_17_retime_s1_44_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_44_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_44_reg_reg_IQ <= mul_34_17_n_10153;
     end
 assign mul_34_17_n_10866 = mul_34_17_retime_s1_44_reg_reg_IQ;
 reg mul_34_17_retime_s1_45_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_45_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_45_reg_reg_IQ <= mul_34_17_n_9984;
     end
 assign mul_34_17_n_10867 = mul_34_17_retime_s1_45_reg_reg_IQ;
 reg mul_34_17_retime_s1_46_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_46_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_46_reg_reg_IQ <= mul_34_17_n_10030;
     end
 assign mul_34_17_n_10868 = mul_34_17_retime_s1_46_reg_reg_IQ;
 reg mul_34_17_retime_s1_47_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_47_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_47_reg_reg_IQ <= mul_34_17_n_10131;
     end
 assign mul_34_17_n_10869 = mul_34_17_retime_s1_47_reg_reg_IQ;
 reg mul_34_17_retime_s1_48_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_48_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_48_reg_reg_IQ <= mul_34_17_n_10137;
     end
 assign mul_34_17_n_10870 = mul_34_17_retime_s1_48_reg_reg_IQ;
 reg mul_34_17_retime_s1_49_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_49_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_49_reg_reg_IQ <= mul_34_17_n_10184;
     end
 assign mul_34_17_n_10871 = mul_34_17_retime_s1_49_reg_reg_IQ;
 reg mul_34_17_retime_s1_50_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_50_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_50_reg_reg_IQ <= mul_34_17_n_10181;
     end
 assign mul_34_17_n_10872 = mul_34_17_retime_s1_50_reg_reg_IQ;
 reg mul_34_17_retime_s1_51_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_51_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_51_reg_reg_IQ <= mul_34_17_n_10226;
     end
 assign mul_34_17_n_10873 = mul_34_17_retime_s1_51_reg_reg_IQ;
 reg mul_34_17_retime_s1_52_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_52_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_52_reg_reg_IQ <= mul_34_17_n_344;
     end
 assign mul_34_17_n_10874 = mul_34_17_retime_s1_52_reg_reg_IQ;
 reg mul_34_17_retime_s1_53_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_53_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_53_reg_reg_IQ <= mul_34_17_n_10094;
     end
 assign mul_34_17_n_10875 = mul_34_17_retime_s1_53_reg_reg_IQ;
 reg mul_34_17_retime_s1_54_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_54_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_54_reg_reg_IQ <= mul_34_17_n_10235;
     end
 assign mul_34_17_n_10876 = mul_34_17_retime_s1_54_reg_reg_IQ;
 reg mul_34_17_retime_s1_55_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_55_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_55_reg_reg_IQ <= mul_34_17_n_10113;
     end
 assign mul_34_17_n_10877 = mul_34_17_retime_s1_55_reg_reg_IQ;
 reg mul_34_17_retime_s1_56_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_56_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_56_reg_reg_IQ <= mul_34_17_n_10152;
     end
 assign mul_34_17_n_10878 = mul_34_17_retime_s1_56_reg_reg_IQ;
 reg mul_34_17_retime_s1_57_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_57_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_57_reg_reg_IQ <= mul_34_17_n_10225;
     end
 assign mul_34_17_n_10879 = mul_34_17_retime_s1_57_reg_reg_IQ;
 reg mul_34_17_retime_s1_58_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_58_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_58_reg_reg_IQ <= mul_34_17_n_10129;
     end
 assign mul_34_17_n_10880 = mul_34_17_retime_s1_58_reg_reg_IQ;
 reg mul_34_17_retime_s1_59_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_59_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_59_reg_reg_IQ <= mul_34_17_n_10257;
     end
 assign mul_34_17_n_10881 = mul_34_17_retime_s1_59_reg_reg_IQ;
 reg mul_34_17_retime_s1_60_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_60_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_60_reg_reg_IQ <= mul_34_17_n_10277;
     end
 assign mul_34_17_n_10882 = mul_34_17_retime_s1_60_reg_reg_IQ;
 reg mul_34_17_retime_s1_61_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_61_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_61_reg_reg_IQ <= mul_34_17_n_10256;
     end
 assign mul_34_17_n_10883 = mul_34_17_retime_s1_61_reg_reg_IQ;
 reg mul_34_17_retime_s1_62_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_62_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_62_reg_reg_IQ <= mul_34_17_n_9951;
     end
 assign mul_34_17_n_10884 = mul_34_17_retime_s1_62_reg_reg_IQ;
 reg mul_34_17_retime_s1_63_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_63_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_63_reg_reg_IQ <= mul_34_17_n_10234;
     end
 assign mul_34_17_n_10885 = mul_34_17_retime_s1_63_reg_reg_IQ;
 reg mul_34_17_retime_s1_64_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_64_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_64_reg_reg_IQ <= mul_34_17_n_10237;
     end
 assign mul_34_17_n_10886 = mul_34_17_retime_s1_64_reg_reg_IQ;
 reg mul_34_17_retime_s1_65_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_65_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_65_reg_reg_IQ <= mul_34_17_n_337;
     end
 assign mul_34_17_n_10887 = mul_34_17_retime_s1_65_reg_reg_IQ;
 reg mul_34_17_retime_s1_66_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_66_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_66_reg_reg_IQ <= mul_34_17_n_10196;
     end
 assign mul_34_17_n_10888 = mul_34_17_retime_s1_66_reg_reg_IQ;
 reg mul_34_17_retime_s1_67_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_67_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_67_reg_reg_IQ <= mul_34_17_n_9865;
     end
 assign mul_34_17_n_10889 = mul_34_17_retime_s1_67_reg_reg_IQ;
 reg mul_34_17_retime_s1_68_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_68_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_68_reg_reg_IQ <= mul_34_17_n_10074;
     end
 assign mul_34_17_n_11252 = mul_34_17_retime_s1_68_reg_reg_IQ;
 reg mul_34_17_retime_s1_69_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_69_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_69_reg_reg_IQ <= mul_34_17_n_10148;
     end
 assign mul_34_17_n_10890 = mul_34_17_retime_s1_69_reg_reg_IQ;
 reg mul_34_17_retime_s1_70_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_70_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_70_reg_reg_IQ <= mul_34_17_n_325;
     end
 assign mul_34_17_n_10891 = mul_34_17_retime_s1_70_reg_reg_IQ;
 reg mul_34_17_retime_s1_71_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_71_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_71_reg_reg_IQ <= mul_34_17_n_10049;
     end
 assign mul_34_17_n_10892 = mul_34_17_retime_s1_71_reg_reg_IQ;
 reg mul_34_17_retime_s1_72_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_72_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_72_reg_reg_IQ <= mul_34_17_n_10263;
     end
 assign mul_34_17_n_10893 = mul_34_17_retime_s1_72_reg_reg_IQ;
 reg mul_34_17_retime_s1_73_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_73_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_73_reg_reg_IQ <= mul_34_17_n_10209;
     end
 assign mul_34_17_n_10894 = mul_34_17_retime_s1_73_reg_reg_IQ;
 reg mul_34_17_retime_s1_74_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_74_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_74_reg_reg_IQ <= mul_34_17_n_10232;
     end
 assign mul_34_17_n_10895 = mul_34_17_retime_s1_74_reg_reg_IQ;
 reg mul_34_17_retime_s1_75_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_75_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_75_reg_reg_IQ <= mul_34_17_n_10262;
     end
 assign mul_34_17_n_10896 = mul_34_17_retime_s1_75_reg_reg_IQ;
 reg mul_34_17_retime_s1_76_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_76_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_76_reg_reg_IQ <= mul_34_17_n_10242;
     end
 assign mul_34_17_n_10897 = mul_34_17_retime_s1_76_reg_reg_IQ;
 reg mul_34_17_retime_s1_77_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_77_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_77_reg_reg_IQ <= mul_34_17_n_10099;
     end
 assign mul_34_17_n_10898 = mul_34_17_retime_s1_77_reg_reg_IQ;
 reg mul_34_17_retime_s1_78_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_78_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_78_reg_reg_IQ <= mul_34_17_n_10239;
     end
 assign mul_34_17_n_10899 = mul_34_17_retime_s1_78_reg_reg_IQ;
 reg mul_34_17_retime_s1_79_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_79_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_79_reg_reg_IQ <= mul_34_17_n_10126;
     end
 assign mul_34_17_n_10900 = mul_34_17_retime_s1_79_reg_reg_IQ;
 reg mul_34_17_retime_s1_80_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_80_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_80_reg_reg_IQ <= mul_34_17_n_10080;
     end
 assign mul_34_17_n_10901 = mul_34_17_retime_s1_80_reg_reg_IQ;
 reg mul_34_17_retime_s1_81_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_81_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_81_reg_reg_IQ <= mul_34_17_n_10045;
     end
 assign mul_34_17_n_10902 = mul_34_17_retime_s1_81_reg_reg_IQ;
 reg mul_34_17_retime_s1_82_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_82_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_82_reg_reg_IQ <= mul_34_17_n_10183;
     end
 assign mul_34_17_n_10903 = mul_34_17_retime_s1_82_reg_reg_IQ;
 reg mul_34_17_retime_s1_83_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_83_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_83_reg_reg_IQ <= mul_34_17_n_10125;
     end
 assign mul_34_17_n_10904 = mul_34_17_retime_s1_83_reg_reg_IQ;
 reg mul_34_17_retime_s1_84_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_84_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_84_reg_reg_IQ <= mul_34_17_n_10182;
     end
 assign mul_34_17_n_10905 = mul_34_17_retime_s1_84_reg_reg_IQ;
 reg mul_34_17_retime_s1_85_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_85_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_85_reg_reg_IQ <= mul_34_17_n_10110;
     end
 assign mul_34_17_n_10906 = mul_34_17_retime_s1_85_reg_reg_IQ;
 reg mul_34_17_retime_s1_86_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_86_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_86_reg_reg_IQ <= mul_34_17_n_9949;
     end
 assign mul_34_17_n_10907 = mul_34_17_retime_s1_86_reg_reg_IQ;
 reg mul_34_17_retime_s1_87_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_87_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_87_reg_reg_IQ <= mul_34_17_n_10180;
     end
 assign mul_34_17_n_10908 = mul_34_17_retime_s1_87_reg_reg_IQ;
 reg mul_34_17_retime_s1_88_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_88_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_88_reg_reg_IQ <= mul_34_17_n_10179;
     end
 assign mul_34_17_n_10909 = mul_34_17_retime_s1_88_reg_reg_IQ;
 reg mul_34_17_retime_s1_89_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_89_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_89_reg_reg_IQ <= mul_34_17_n_10203;
     end
 assign mul_34_17_n_10910 = mul_34_17_retime_s1_89_reg_reg_IQ;
 reg mul_34_17_retime_s1_90_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_90_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_90_reg_reg_IQ <= mul_34_17_n_10208;
     end
 assign mul_34_17_n_10911 = mul_34_17_retime_s1_90_reg_reg_IQ;
 reg mul_34_17_retime_s1_91_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_91_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_91_reg_reg_IQ <= mul_34_17_n_10276;
     end
 assign mul_34_17_n_10912 = mul_34_17_retime_s1_91_reg_reg_IQ;
 reg mul_34_17_retime_s1_92_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_92_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_92_reg_reg_IQ <= mul_34_17_n_10216;
     end
 assign mul_34_17_n_10913 = mul_34_17_retime_s1_92_reg_reg_IQ;
 reg mul_34_17_retime_s1_93_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_93_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_93_reg_reg_IQ <= mul_34_17_n_10275;
     end
 assign mul_34_17_n_10914 = mul_34_17_retime_s1_93_reg_reg_IQ;
 reg mul_34_17_retime_s1_94_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_94_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_94_reg_reg_IQ <= mul_34_17_n_10252;
     end
 assign mul_34_17_n_10915 = mul_34_17_retime_s1_94_reg_reg_IQ;
 reg mul_34_17_retime_s1_95_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_95_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_95_reg_reg_IQ <= mul_34_17_n_10146;
     end
 assign mul_34_17_n_10916 = mul_34_17_retime_s1_95_reg_reg_IQ;
 reg mul_34_17_retime_s1_96_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_96_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_96_reg_reg_IQ <= mul_34_17_n_10022;
     end
 assign mul_34_17_n_10917 = mul_34_17_retime_s1_96_reg_reg_IQ;
 reg mul_34_17_retime_s1_97_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_97_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_97_reg_reg_IQ <= mul_34_17_n_10195;
     end
 assign mul_34_17_n_10918 = mul_34_17_retime_s1_97_reg_reg_IQ;
 reg mul_34_17_retime_s1_98_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_98_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_98_reg_reg_IQ <= mul_34_17_n_10145;
     end
 assign mul_34_17_n_10919 = mul_34_17_retime_s1_98_reg_reg_IQ;
 reg mul_34_17_retime_s1_99_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_99_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_99_reg_reg_IQ <= mul_34_17_n_10164;
     end
 assign mul_34_17_n_10920 = mul_34_17_retime_s1_99_reg_reg_IQ;
 reg mul_34_17_retime_s1_100_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_100_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_100_reg_reg_IQ <= mul_34_17_n_9988;
     end
 assign mul_34_17_n_11253 = mul_34_17_retime_s1_100_reg_reg_IQ;
 reg mul_34_17_retime_s1_101_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_101_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_101_reg_reg_IQ <= mul_34_17_n_10069;
     end
 assign mul_34_17_n_10921 = mul_34_17_retime_s1_101_reg_reg_IQ;
 reg mul_34_17_retime_s1_102_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_102_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_102_reg_reg_IQ <= mul_34_17_n_10273;
     end
 assign mul_34_17_n_10922 = mul_34_17_retime_s1_102_reg_reg_IQ;
 reg mul_34_17_retime_s1_103_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_103_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_103_reg_reg_IQ <= mul_34_17_n_10255;
     end
 assign mul_34_17_n_10923 = mul_34_17_retime_s1_103_reg_reg_IQ;
 reg mul_34_17_retime_s1_104_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_104_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_104_reg_reg_IQ <= mul_34_17_n_10274;
     end
 assign mul_34_17_n_10924 = mul_34_17_retime_s1_104_reg_reg_IQ;
 reg mul_34_17_retime_s1_105_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_105_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_105_reg_reg_IQ <= mul_34_17_n_10243;
     end
 assign mul_34_17_n_10925 = mul_34_17_retime_s1_105_reg_reg_IQ;
 reg mul_34_17_retime_s1_106_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_106_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_106_reg_reg_IQ <= mul_34_17_n_9677;
     end
 assign mul_34_17_n_10926 = mul_34_17_retime_s1_106_reg_reg_IQ;
 reg mul_34_17_retime_s1_107_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_107_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_107_reg_reg_IQ <= mul_34_17_n_9518;
     end
 assign mul_34_17_n_10927 = mul_34_17_retime_s1_107_reg_reg_IQ;
 reg mul_34_17_retime_s1_108_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_108_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_108_reg_reg_IQ <= mul_34_17_n_10090;
     end
 assign mul_34_17_n_10928 = mul_34_17_retime_s1_108_reg_reg_IQ;
 reg mul_34_17_retime_s1_109_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_109_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_109_reg_reg_IQ <= mul_34_17_n_10177;
     end
 assign mul_34_17_n_10929 = mul_34_17_retime_s1_109_reg_reg_IQ;
 reg mul_34_17_retime_s1_110_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_110_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_110_reg_reg_IQ <= mul_34_17_n_10178;
     end
 assign mul_34_17_n_10930 = mul_34_17_retime_s1_110_reg_reg_IQ;
 reg mul_34_17_retime_s1_111_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_111_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_111_reg_reg_IQ <= mul_34_17_n_10073;
     end
 assign mul_34_17_n_10931 = mul_34_17_retime_s1_111_reg_reg_IQ;
 reg mul_34_17_retime_s1_112_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_112_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_112_reg_reg_IQ <= mul_34_17_n_9683;
     end
 assign mul_34_17_n_10932 = mul_34_17_retime_s1_112_reg_reg_IQ;
 reg mul_34_17_retime_s1_113_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_113_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_113_reg_reg_IQ <= mul_34_17_n_9934;
     end
 assign mul_34_17_n_10933 = mul_34_17_retime_s1_113_reg_reg_IQ;
 reg mul_34_17_retime_s1_114_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_114_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_114_reg_reg_IQ <= mul_34_17_n_9989;
     end
 assign mul_34_17_n_10934 = mul_34_17_retime_s1_114_reg_reg_IQ;
 reg mul_34_17_retime_s1_115_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_115_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_115_reg_reg_IQ <= mul_34_17_n_9963;
     end
 assign mul_34_17_n_10935 = mul_34_17_retime_s1_115_reg_reg_IQ;
 reg mul_34_17_retime_s1_116_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_116_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_116_reg_reg_IQ <= mul_34_17_n_10043;
     end
 assign mul_34_17_n_10936 = mul_34_17_retime_s1_116_reg_reg_IQ;
 reg mul_34_17_retime_s1_117_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_117_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_117_reg_reg_IQ <= mul_34_17_n_9623;
     end
 assign mul_34_17_n_10937 = mul_34_17_retime_s1_117_reg_reg_IQ;
 reg mul_34_17_retime_s1_118_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_118_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_118_reg_reg_IQ <= mul_34_17_n_9607;
     end
 assign mul_34_17_n_10938 = mul_34_17_retime_s1_118_reg_reg_IQ;
 reg mul_34_17_retime_s1_119_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_119_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_119_reg_reg_IQ <= mul_34_17_n_10202;
     end
 assign mul_34_17_n_10939 = mul_34_17_retime_s1_119_reg_reg_IQ;
 reg mul_34_17_retime_s1_120_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_120_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_120_reg_reg_IQ <= mul_34_17_n_10261;
     end
 assign mul_34_17_n_10940 = mul_34_17_retime_s1_120_reg_reg_IQ;
 reg mul_34_17_retime_s1_121_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_121_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_121_reg_reg_IQ <= mul_34_17_n_10201;
     end
 assign mul_34_17_n_10941 = mul_34_17_retime_s1_121_reg_reg_IQ;
 reg mul_34_17_retime_s1_122_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_122_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_122_reg_reg_IQ <= mul_34_17_n_10272;
     end
 assign mul_34_17_n_10942 = mul_34_17_retime_s1_122_reg_reg_IQ;
 reg mul_34_17_retime_s1_123_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_123_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_123_reg_reg_IQ <= mul_34_17_n_2872;
     end
 assign mul_34_17_n_10943 = mul_34_17_retime_s1_123_reg_reg_IQ;
 reg mul_34_17_retime_s1_124_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_124_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_124_reg_reg_IQ <= mul_34_17_n_10260;
     end
 assign mul_34_17_n_10944 = mul_34_17_retime_s1_124_reg_reg_IQ;
 reg mul_34_17_retime_s1_125_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_125_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_125_reg_reg_IQ <= mul_34_17_n_10105;
     end
 assign mul_34_17_n_10945 = mul_34_17_retime_s1_125_reg_reg_IQ;
 reg mul_34_17_retime_s1_126_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_126_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_126_reg_reg_IQ <= mul_34_17_n_10222;
     end
 assign mul_34_17_n_10946 = mul_34_17_retime_s1_126_reg_reg_IQ;
 reg mul_34_17_retime_s1_127_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_127_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_127_reg_reg_IQ <= mul_34_17_n_10143;
     end
 assign mul_34_17_n_10947 = mul_34_17_retime_s1_127_reg_reg_IQ;
 reg mul_34_17_retime_s1_128_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_128_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_128_reg_reg_IQ <= mul_34_17_n_10151;
     end
 assign mul_34_17_n_10948 = mul_34_17_retime_s1_128_reg_reg_IQ;
 reg mul_34_17_retime_s1_129_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_129_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_129_reg_reg_IQ <= mul_34_17_n_10200;
     end
 assign mul_34_17_n_10949 = mul_34_17_retime_s1_129_reg_reg_IQ;
 reg mul_34_17_retime_s1_130_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_130_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_130_reg_reg_IQ <= mul_34_17_n_339;
     end
 assign mul_34_17_n_10950 = mul_34_17_retime_s1_130_reg_reg_IQ;
 reg mul_34_17_retime_s1_131_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_131_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_131_reg_reg_IQ <= mul_34_17_n_10199;
     end
 assign mul_34_17_n_10951 = mul_34_17_retime_s1_131_reg_reg_IQ;
 reg mul_34_17_retime_s1_132_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_132_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_132_reg_reg_IQ <= mul_34_17_n_327;
     end
 assign mul_34_17_n_10952 = mul_34_17_retime_s1_132_reg_reg_IQ;
 reg mul_34_17_retime_s1_133_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_133_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_133_reg_reg_IQ <= mul_34_17_n_10155;
     end
 assign mul_34_17_n_10953 = mul_34_17_retime_s1_133_reg_reg_IQ;
 reg mul_34_17_retime_s1_134_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_134_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_134_reg_reg_IQ <= mul_34_17_n_9914;
     end
 assign mul_34_17_n_10954 = mul_34_17_retime_s1_134_reg_reg_IQ;
 reg mul_34_17_retime_s1_135_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_135_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_135_reg_reg_IQ <= mul_34_17_n_328;
     end
 assign mul_34_17_n_10955 = mul_34_17_retime_s1_135_reg_reg_IQ;
 reg mul_34_17_retime_s1_136_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_136_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_136_reg_reg_IQ <= mul_34_17_n_9857;
     end
 assign mul_34_17_n_10956 = mul_34_17_retime_s1_136_reg_reg_IQ;
 reg mul_34_17_retime_s1_137_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_137_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_137_reg_reg_IQ <= mul_34_17_n_9964;
     end
 assign mul_34_17_n_10957 = mul_34_17_retime_s1_137_reg_reg_IQ;
 reg mul_34_17_retime_s1_138_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_138_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_138_reg_reg_IQ <= mul_34_17_n_9362;
     end
 assign mul_34_17_n_10958 = mul_34_17_retime_s1_138_reg_reg_IQ;
 reg mul_34_17_retime_s1_139_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_139_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_139_reg_reg_IQ <= mul_34_17_n_9543;
     end
 assign mul_34_17_n_10959 = mul_34_17_retime_s1_139_reg_reg_IQ;
 reg mul_34_17_retime_s1_140_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_140_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_140_reg_reg_IQ <= mul_34_17_n_9652;
     end
 assign mul_34_17_n_10960 = mul_34_17_retime_s1_140_reg_reg_IQ;
 reg mul_34_17_retime_s1_141_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_141_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_141_reg_reg_IQ <= mul_34_17_n_9645;
     end
 assign mul_34_17_n_10961 = mul_34_17_retime_s1_141_reg_reg_IQ;
 reg mul_34_17_retime_s1_142_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_142_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_142_reg_reg_IQ <= mul_34_17_n_9438;
     end
 assign mul_34_17_n_10962 = mul_34_17_retime_s1_142_reg_reg_IQ;
 reg mul_34_17_retime_s1_143_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_143_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_143_reg_reg_IQ <= mul_34_17_n_9751;
     end
 assign mul_34_17_n_10963 = mul_34_17_retime_s1_143_reg_reg_IQ;
 reg mul_34_17_retime_s1_144_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_144_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_144_reg_reg_IQ <= mul_34_17_n_10221;
     end
 assign mul_34_17_n_10964 = mul_34_17_retime_s1_144_reg_reg_IQ;
 reg mul_34_17_retime_s1_145_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_145_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_145_reg_reg_IQ <= mul_34_17_n_9704;
     end
 assign mul_34_17_n_10965 = mul_34_17_retime_s1_145_reg_reg_IQ;
 reg mul_34_17_retime_s1_146_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_146_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_146_reg_reg_IQ <= mul_34_17_n_9456;
     end
 assign mul_34_17_n_10966 = mul_34_17_retime_s1_146_reg_reg_IQ;
 reg mul_34_17_retime_s1_147_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_147_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_147_reg_reg_IQ <= mul_34_17_n_9942;
     end
 assign mul_34_17_n_10967 = mul_34_17_retime_s1_147_reg_reg_IQ;
 reg mul_34_17_retime_s1_148_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_148_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_148_reg_reg_IQ <= mul_34_17_n_9941;
     end
 assign mul_34_17_n_10968 = mul_34_17_retime_s1_148_reg_reg_IQ;
 reg mul_34_17_retime_s1_149_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_149_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_149_reg_reg_IQ <= mul_34_17_n_9972;
     end
 assign mul_34_17_n_10969 = mul_34_17_retime_s1_149_reg_reg_IQ;
 reg mul_34_17_retime_s1_150_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_150_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_150_reg_reg_IQ <= mul_34_17_n_9848;
     end
 assign mul_34_17_n_10970 = mul_34_17_retime_s1_150_reg_reg_IQ;
 reg mul_34_17_retime_s1_151_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_151_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_151_reg_reg_IQ <= mul_34_17_n_10040;
     end
 assign mul_34_17_n_10971 = mul_34_17_retime_s1_151_reg_reg_IQ;
 reg mul_34_17_retime_s1_152_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_152_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_152_reg_reg_IQ <= mul_34_17_n_10053;
     end
 assign mul_34_17_n_10972 = mul_34_17_retime_s1_152_reg_reg_IQ;
 reg mul_34_17_retime_s1_153_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_153_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_153_reg_reg_IQ <= mul_34_17_n_10079;
     end
 assign mul_34_17_n_11251 = mul_34_17_retime_s1_153_reg_reg_IQ;
 reg mul_34_17_retime_s1_154_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_154_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_154_reg_reg_IQ <= mul_34_17_n_9750;
     end
 assign mul_34_17_n_10973 = mul_34_17_retime_s1_154_reg_reg_IQ;
 reg mul_34_17_retime_s1_155_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_155_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_155_reg_reg_IQ <= mul_34_17_n_8279;
     end
 assign mul_34_17_n_10974 = mul_34_17_retime_s1_155_reg_reg_IQ;
 reg mul_34_17_retime_s1_156_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_156_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_156_reg_reg_IQ <= mul_34_17_n_8699;
     end
 assign mul_34_17_n_10975 = mul_34_17_retime_s1_156_reg_reg_IQ;
 reg mul_34_17_retime_s1_157_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_157_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_157_reg_reg_IQ <= mul_34_17_n_8798;
     end
 assign mul_34_17_n_10976 = mul_34_17_retime_s1_157_reg_reg_IQ;
 reg mul_34_17_retime_s1_158_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_158_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_158_reg_reg_IQ <= mul_34_17_n_9302;
     end
 assign mul_34_17_n_10977 = mul_34_17_retime_s1_158_reg_reg_IQ;
 reg mul_34_17_retime_s1_159_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_159_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_159_reg_reg_IQ <= mul_34_17_n_9073;
     end
 assign mul_34_17_n_10978 = mul_34_17_retime_s1_159_reg_reg_IQ;
 reg mul_34_17_retime_s1_160_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_160_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_160_reg_reg_IQ <= mul_34_17_n_9072;
     end
 assign mul_34_17_n_10979 = mul_34_17_retime_s1_160_reg_reg_IQ;
 reg mul_34_17_retime_s1_161_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_161_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_161_reg_reg_IQ <= mul_34_17_n_9753;
     end
 assign mul_34_17_n_10980 = mul_34_17_retime_s1_161_reg_reg_IQ;
 reg mul_34_17_retime_s1_162_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_162_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_162_reg_reg_IQ <= mul_34_17_n_9212;
     end
 assign mul_34_17_n_10981 = mul_34_17_retime_s1_162_reg_reg_IQ;
 reg mul_34_17_retime_s1_163_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_163_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_163_reg_reg_IQ <= mul_34_17_n_9153;
     end
 assign mul_34_17_n_10982 = mul_34_17_retime_s1_163_reg_reg_IQ;
 reg mul_34_17_retime_s1_164_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_164_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_164_reg_reg_IQ <= mul_34_17_n_10122;
     end
 assign mul_34_17_n_10983 = mul_34_17_retime_s1_164_reg_reg_IQ;
 reg mul_34_17_retime_s1_165_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_165_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_165_reg_reg_IQ <= mul_34_17_n_9079;
     end
 assign mul_34_17_n_10984 = mul_34_17_retime_s1_165_reg_reg_IQ;
 reg mul_34_17_retime_s1_166_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_166_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_166_reg_reg_IQ <= mul_34_17_n_8308;
     end
 assign mul_34_17_n_10985 = mul_34_17_retime_s1_166_reg_reg_IQ;
 reg mul_34_17_retime_s1_167_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_167_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_167_reg_reg_IQ <= mul_34_17_n_7274;
     end
 assign mul_34_17_n_10986 = mul_34_17_retime_s1_167_reg_reg_IQ;
 reg mul_34_17_retime_s1_168_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_168_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_168_reg_reg_IQ <= mul_34_17_n_7624;
     end
 assign mul_34_17_n_10987 = mul_34_17_retime_s1_168_reg_reg_IQ;
 reg mul_34_17_retime_s1_169_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_169_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_169_reg_reg_IQ <= mul_34_17_n_518;
     end
 assign asc001_0_ = mul_34_17_retime_s1_169_reg_reg_IQ;
 reg mul_34_17_retime_s1_170_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_170_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_170_reg_reg_IQ <= mul_34_17_n_2239;
     end
 assign mul_34_17_n_10988 = mul_34_17_retime_s1_170_reg_reg_IQ;
 reg mul_34_17_retime_s1_171_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_171_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_171_reg_reg_IQ <= mul_34_17_n_9259;
     end
 assign mul_34_17_n_10989 = mul_34_17_retime_s1_171_reg_reg_IQ;
 reg mul_34_17_retime_s1_172_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_172_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_172_reg_reg_IQ <= mul_34_17_n_9249;
     end
 assign mul_34_17_n_10990 = mul_34_17_retime_s1_172_reg_reg_IQ;
 reg mul_34_17_retime_s1_173_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_173_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_173_reg_reg_IQ <= mul_34_17_n_9939;
     end
 assign mul_34_17_n_10991 = mul_34_17_retime_s1_173_reg_reg_IQ;
 reg mul_34_17_retime_s1_174_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_174_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_174_reg_reg_IQ <= mul_34_17_n_321;
     end
 assign mul_34_17_n_10992 = mul_34_17_retime_s1_174_reg_reg_IQ;
 reg mul_34_17_retime_s1_175_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_175_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_175_reg_reg_IQ <= mul_34_17_n_9938;
     end
 assign mul_34_17_n_10993 = mul_34_17_retime_s1_175_reg_reg_IQ;
 reg mul_34_17_retime_s1_176_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_176_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_176_reg_reg_IQ <= mul_34_17_n_10268;
     end
 assign mul_34_17_n_10994 = mul_34_17_retime_s1_176_reg_reg_IQ;
 reg mul_34_17_retime_s1_177_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_177_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_177_reg_reg_IQ <= mul_34_17_n_10150;
     end
 assign mul_34_17_n_10995 = mul_34_17_retime_s1_177_reg_reg_IQ;
 reg mul_34_17_retime_s1_178_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_178_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_178_reg_reg_IQ <= mul_34_17_n_10020;
     end
 assign mul_34_17_n_10996 = mul_34_17_retime_s1_178_reg_reg_IQ;
 reg mul_34_17_retime_s1_179_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_179_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_179_reg_reg_IQ <= mul_34_17_n_10121;
     end
 assign mul_34_17_n_10997 = mul_34_17_retime_s1_179_reg_reg_IQ;
 reg mul_34_17_retime_s1_180_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_180_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_180_reg_reg_IQ <= mul_34_17_n_10231;
     end
 assign mul_34_17_n_10998 = mul_34_17_retime_s1_180_reg_reg_IQ;
 reg mul_34_17_retime_s1_181_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_181_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_181_reg_reg_IQ <= mul_34_17_n_10120;
     end
 assign mul_34_17_n_10999 = mul_34_17_retime_s1_181_reg_reg_IQ;
 reg mul_34_17_retime_s1_182_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_182_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_182_reg_reg_IQ <= mul_34_17_n_9808;
     end
 assign mul_34_17_n_11000 = mul_34_17_retime_s1_182_reg_reg_IQ;
 reg mul_34_17_retime_s1_183_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_183_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_183_reg_reg_IQ <= mul_34_17_n_10161;
     end
 assign mul_34_17_n_11001 = mul_34_17_retime_s1_183_reg_reg_IQ;
 reg mul_34_17_retime_s1_184_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_184_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_184_reg_reg_IQ <= mul_34_17_n_10037;
     end
 assign mul_34_17_n_11002 = mul_34_17_retime_s1_184_reg_reg_IQ;
 reg mul_34_17_retime_s1_185_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_185_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_185_reg_reg_IQ <= mul_34_17_n_335;
     end
 assign mul_34_17_n_11003 = mul_34_17_retime_s1_185_reg_reg_IQ;
 reg mul_34_17_retime_s1_186_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_186_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_186_reg_reg_IQ <= mul_34_17_n_10267;
     end
 assign mul_34_17_n_11004 = mul_34_17_retime_s1_186_reg_reg_IQ;
 reg mul_34_17_retime_s1_187_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_187_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_187_reg_reg_IQ <= mul_34_17_n_10038;
     end
 assign mul_34_17_n_11005 = mul_34_17_retime_s1_187_reg_reg_IQ;
 reg mul_34_17_retime_s1_188_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_188_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_188_reg_reg_IQ <= mul_34_17_n_9987;
     end
 assign mul_34_17_n_11006 = mul_34_17_retime_s1_188_reg_reg_IQ;
 reg mul_34_17_retime_s1_189_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_189_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_189_reg_reg_IQ <= mul_34_17_n_10198;
     end
 assign mul_34_17_n_11007 = mul_34_17_retime_s1_189_reg_reg_IQ;
 reg mul_34_17_retime_s1_190_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_190_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_190_reg_reg_IQ <= mul_34_17_n_10170;
     end
 assign mul_34_17_n_11008 = mul_34_17_retime_s1_190_reg_reg_IQ;
 reg mul_34_17_retime_s1_191_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_191_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_191_reg_reg_IQ <= mul_34_17_n_9525;
     end
 assign mul_34_17_n_11009 = mul_34_17_retime_s1_191_reg_reg_IQ;
 reg mul_34_17_retime_s1_192_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_192_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_192_reg_reg_IQ <= mul_34_17_n_8470;
     end
 assign mul_34_17_n_11010 = mul_34_17_retime_s1_192_reg_reg_IQ;
 reg mul_34_17_retime_s1_193_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_193_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_193_reg_reg_IQ <= mul_34_17_n_10119;
     end
 assign mul_34_17_n_11011 = mul_34_17_retime_s1_193_reg_reg_IQ;
 reg mul_34_17_retime_s1_194_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_194_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_194_reg_reg_IQ <= mul_34_17_n_7975;
     end
 assign mul_34_17_n_11012 = mul_34_17_retime_s1_194_reg_reg_IQ;
 reg mul_34_17_retime_s1_195_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_195_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_195_reg_reg_IQ <= mul_34_17_n_3039;
     end
 assign mul_34_17_n_11013 = mul_34_17_retime_s1_195_reg_reg_IQ;
 reg mul_34_17_retime_s1_196_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_196_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_196_reg_reg_IQ <= mul_34_17_n_9754;
     end
 assign mul_34_17_n_11014 = mul_34_17_retime_s1_196_reg_reg_IQ;
 reg mul_34_17_retime_s1_197_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_197_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_197_reg_reg_IQ <= mul_34_17_n_9494;
     end
 assign mul_34_17_n_11015 = mul_34_17_retime_s1_197_reg_reg_IQ;
 reg mul_34_17_retime_s1_198_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_198_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_198_reg_reg_IQ <= mul_34_17_n_10204;
     end
 assign mul_34_17_n_11016 = mul_34_17_retime_s1_198_reg_reg_IQ;
 reg mul_34_17_retime_s1_199_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_199_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_199_reg_reg_IQ <= mul_34_17_n_10147;
     end
 assign mul_34_17_n_11017 = mul_34_17_retime_s1_199_reg_reg_IQ;
 reg mul_34_17_retime_s1_200_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_200_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_200_reg_reg_IQ <= mul_34_17_n_9856;
     end
 assign mul_34_17_n_11018 = mul_34_17_retime_s1_200_reg_reg_IQ;
 reg mul_34_17_retime_s1_201_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_201_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_201_reg_reg_IQ <= mul_34_17_n_10165;
     end
 assign mul_34_17_n_11019 = mul_34_17_retime_s1_201_reg_reg_IQ;
 reg mul_34_17_retime_s1_202_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_202_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_202_reg_reg_IQ <= mul_34_17_n_10149;
     end
 assign mul_34_17_n_11020 = mul_34_17_retime_s1_202_reg_reg_IQ;
 reg mul_34_17_retime_s1_203_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_203_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_203_reg_reg_IQ <= mul_34_17_n_10211;
     end
 assign mul_34_17_n_11021 = mul_34_17_retime_s1_203_reg_reg_IQ;
 reg mul_34_17_retime_s1_204_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_204_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_204_reg_reg_IQ <= mul_34_17_n_10266;
     end
 assign mul_34_17_n_11022 = mul_34_17_retime_s1_204_reg_reg_IQ;
 reg mul_34_17_retime_s1_205_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_205_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_205_reg_reg_IQ <= mul_34_17_n_10213;
     end
 assign mul_34_17_n_11023 = mul_34_17_retime_s1_205_reg_reg_IQ;
 reg mul_34_17_retime_s1_206_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_206_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_206_reg_reg_IQ <= mul_34_17_n_10279;
     end
 assign mul_34_17_n_11024 = mul_34_17_retime_s1_206_reg_reg_IQ;
 reg mul_34_17_retime_s1_207_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_207_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_207_reg_reg_IQ <= mul_34_17_n_10212;
     end
 assign mul_34_17_n_11025 = mul_34_17_retime_s1_207_reg_reg_IQ;
 reg mul_34_17_retime_s1_208_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_208_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_208_reg_reg_IQ <= mul_34_17_n_7974;
     end
 assign mul_34_17_n_11026 = mul_34_17_retime_s1_208_reg_reg_IQ;
 reg mul_34_17_retime_s1_209_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_209_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_209_reg_reg_IQ <= mul_34_17_n_7253;
     end
 assign mul_34_17_n_11027 = mul_34_17_retime_s1_209_reg_reg_IQ;
 reg mul_34_17_retime_s1_210_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_210_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_210_reg_reg_IQ <= mul_34_17_n_10117;
     end
 assign mul_34_17_n_11028 = mul_34_17_retime_s1_210_reg_reg_IQ;
 reg mul_34_17_retime_s1_211_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_211_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_211_reg_reg_IQ <= mul_34_17_n_10118;
     end
 assign mul_34_17_n_11029 = mul_34_17_retime_s1_211_reg_reg_IQ;
 reg mul_34_17_retime_s1_212_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_212_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_212_reg_reg_IQ <= mul_34_17_n_330;
     end
 assign mul_34_17_n_11030 = mul_34_17_retime_s1_212_reg_reg_IQ;
 reg mul_34_17_retime_s1_213_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_213_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_213_reg_reg_IQ <= mul_34_17_n_346;
     end
 assign mul_34_17_n_11031 = mul_34_17_retime_s1_213_reg_reg_IQ;
 reg mul_34_17_retime_s1_214_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_214_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_214_reg_reg_IQ <= mul_34_17_n_10223;
     end
 assign mul_34_17_n_11032 = mul_34_17_retime_s1_214_reg_reg_IQ;
 reg mul_34_17_retime_s1_215_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_215_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_215_reg_reg_IQ <= mul_34_17_n_10233;
     end
 assign mul_34_17_n_11033 = mul_34_17_retime_s1_215_reg_reg_IQ;
 reg mul_34_17_retime_s1_216_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_216_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_216_reg_reg_IQ <= mul_34_17_n_10127;
     end
 assign mul_34_17_n_11034 = mul_34_17_retime_s1_216_reg_reg_IQ;
 reg mul_34_17_retime_s1_217_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_217_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_217_reg_reg_IQ <= mul_34_17_n_10186;
     end
 assign mul_34_17_n_11035 = mul_34_17_retime_s1_217_reg_reg_IQ;
 reg mul_34_17_retime_s1_218_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_218_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_218_reg_reg_IQ <= mul_34_17_n_303;
     end
 assign mul_34_17_n_11036 = mul_34_17_retime_s1_218_reg_reg_IQ;
 reg mul_34_17_retime_s1_219_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_219_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_219_reg_reg_IQ <= mul_34_17_n_3959;
     end
 assign mul_34_17_n_11037 = mul_34_17_retime_s1_219_reg_reg_IQ;
 reg mul_34_17_retime_s1_220_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_220_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_220_reg_reg_IQ <= mul_34_17_n_10241;
     end
 assign mul_34_17_n_11038 = mul_34_17_retime_s1_220_reg_reg_IQ;
 reg mul_34_17_retime_s1_221_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_221_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_221_reg_reg_IQ <= mul_34_17_n_7384;
     end
 assign mul_34_17_n_11039 = mul_34_17_retime_s1_221_reg_reg_IQ;
 reg mul_34_17_retime_s1_222_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_222_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_222_reg_reg_IQ <= mul_34_17_n_6875;
     end
 assign mul_34_17_n_11040 = mul_34_17_retime_s1_222_reg_reg_IQ;
 reg mul_34_17_retime_s1_223_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_223_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_223_reg_reg_IQ <= mul_34_17_n_10265;
     end
 assign mul_34_17_n_11041 = mul_34_17_retime_s1_223_reg_reg_IQ;
 reg mul_34_17_retime_s1_224_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_224_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_224_reg_reg_IQ <= mul_34_17_n_10116;
     end
 assign mul_34_17_n_11042 = mul_34_17_retime_s1_224_reg_reg_IQ;
 reg mul_34_17_retime_s1_225_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_225_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_225_reg_reg_IQ <= mul_34_17_n_10271;
     end
 assign mul_34_17_n_11043 = mul_34_17_retime_s1_225_reg_reg_IQ;
 reg mul_34_17_retime_s1_226_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_226_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_226_reg_reg_IQ <= mul_34_17_n_10032;
     end
 assign mul_34_17_n_11044 = mul_34_17_retime_s1_226_reg_reg_IQ;
 reg mul_34_17_retime_s1_227_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_227_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_227_reg_reg_IQ <= mul_34_17_n_9762;
     end
 assign mul_34_17_n_11045 = mul_34_17_retime_s1_227_reg_reg_IQ;
 reg mul_34_17_retime_s1_228_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_228_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_228_reg_reg_IQ <= mul_34_17_n_10264;
     end
 assign mul_34_17_n_11046 = mul_34_17_retime_s1_228_reg_reg_IQ;
 reg mul_34_17_retime_s1_229_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_229_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_229_reg_reg_IQ <= mul_34_17_n_10197;
     end
 assign mul_34_17_n_11047 = mul_34_17_retime_s1_229_reg_reg_IQ;
 reg mul_34_17_retime_s1_230_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_230_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_230_reg_reg_IQ <= mul_34_17_n_4875;
     end
 assign mul_34_17_n_11048 = mul_34_17_retime_s1_230_reg_reg_IQ;
 reg mul_34_17_retime_s1_231_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_231_reg_reg_IQ <= 1'B0;
     else begin
         mul_34_17_retime_s1_231_reg_reg_IQ <= mul_34_17_n_10210;
     end
 assign mul_34_17_n_11049 = mul_34_17_retime_s1_231_reg_reg_IQ;
 reg mul_34_17_retime_s1_232_reg_reg_IQ;
 always @(posedge clk or negedge clr)
     if (clr == 1'B0) mul_34_17_retime_s1_232_reg_reg_IQ <= 1'B1;
     else begin
         mul_34_17_retime_s1_232_reg_reg_IQ <= mul_34_17_n_348;
     end
 assign mul_34_17_n_11050 = mul_34_17_retime_s1_232_reg_reg_IQ;
 assign asc001_85_ = (mul_34_17_n_10822 ^ mul_34_17_n_10853);
 assign asc001_75_ = ~(mul_34_17_n_10824 ^ mul_34_17_n_10455);
 assign asc001_84_ = ~(mul_34_17_n_10823 ^ mul_34_17_n_10425);
 assign asc001_83_ = ~(mul_34_17_n_10821 ^ mul_34_17_n_10445);
 assign asc001_82_ = ~(mul_34_17_n_10820 ^ mul_34_17_n_10546);
 assign asc001_81_ = ~(mul_34_17_n_10819 ^ mul_34_17_n_10432);
 assign asc001_74_ = ~(mul_34_17_n_10815 ^ mul_34_17_n_10461);
 assign asc001_76_ = ~(mul_34_17_n_10814 ^ mul_34_17_n_10329);
 assign asc001_77_ = ~(mul_34_17_n_10813 ^ mul_34_17_n_10334);
 assign asc001_73_ = ~(mul_34_17_n_10807 ^ mul_34_17_n_10453);
 assign asc001_69_ = ~(mul_34_17_n_10808 ^ mul_34_17_n_10566);
 assign asc001_70_ = ~(mul_34_17_n_10806 ^ mul_34_17_n_10451);
 assign asc001_71_ = ~(mul_34_17_n_10816 ^ mul_34_17_n_10497);
 assign asc001_79_ = ~(mul_34_17_n_10812 ^ mul_34_17_n_10544);
 assign mul_34_17_n_10824 = ~(mul_34_17_n_10817 & mul_34_17_n_10631);
 assign mul_34_17_n_10823 = ~(mul_34_17_n_10818 & mul_34_17_n_10667);
 assign mul_34_17_n_10822 = ~(mul_34_17_n_10810 & mul_34_17_n_10803);
 assign mul_34_17_n_10821 = ~(mul_34_17_n_10811 & mul_34_17_n_10796);
 assign mul_34_17_n_10820 = ~(mul_34_17_n_10809 & mul_34_17_n_10591);
 assign mul_34_17_n_10819 = ((mul_34_17_n_10435 & mul_34_17_n_10804) | ((mul_34_17_n_10435 & mul_34_17_n_10362)
    | (mul_34_17_n_10362 & mul_34_17_n_10804)));
 assign asc001_78_ = ~(mul_34_17_n_10798 ^ mul_34_17_n_10431);
 assign asc001_63_ = ~(mul_34_17_n_10793 ^ mul_34_17_n_10449);
 assign asc001_62_ = ~(mul_34_17_n_10792 ^ mul_34_17_n_10448);
 assign asc001_61_ = ~(mul_34_17_n_10800 ^ mul_34_17_n_10442);
 assign asc001_59_ = ~(mul_34_17_n_10801 ^ mul_34_17_n_10496);
 assign asc001_80_ = ~(mul_34_17_n_10804 ^ mul_34_17_n_10545);
 assign asc001_67_ = ~(mul_34_17_n_10799 ^ mul_34_17_n_10620);
 assign mul_34_17_n_10818 = ~(mul_34_17_n_10804 & mul_34_17_n_10598);
 assign mul_34_17_n_10817 = ~(mul_34_17_n_10805 & mul_34_17_n_10380);
 assign mul_34_17_n_10816 = ~(mul_34_17_n_10797 | mul_34_17_n_10712);
 assign mul_34_17_n_10815 = ~(mul_34_17_n_10805 | mul_34_17_n_10562);
 assign mul_34_17_n_10814 = ~(mul_34_17_n_10802 | mul_34_17_n_10671);
 assign mul_34_17_n_10813 = ~(mul_34_17_n_10794 | mul_34_17_n_10773);
 assign mul_34_17_n_10812 = ~(mul_34_17_n_10684 | (mul_34_17_n_10500 | (mul_34_17_n_10353 | mul_34_17_n_10795)));
 assign mul_34_17_n_10811 = ((mul_34_17_n_10591 | mul_34_17_n_10528) & (mul_34_17_n_10791 | mul_34_17_n_10610));
 assign mul_34_17_n_10810 = ((mul_34_17_n_10667 | mul_34_17_n_11247) & (mul_34_17_n_10791 | mul_34_17_n_10647));
 assign asc001_72_ = ~(mul_34_17_n_10789 ^ mul_34_17_n_10498);
 assign mul_34_17_n_10809 = ~(mul_34_17_n_10804 & mul_34_17_n_10575);
 assign mul_34_17_n_10808 = ((mul_34_17_n_10511 & mul_34_17_n_10790) | ((mul_34_17_n_10511 & mul_34_17_n_10436)
    | (mul_34_17_n_10436 & mul_34_17_n_10790)));
 assign mul_34_17_n_10807 = ((mul_34_17_n_10400 | mul_34_17_n_10404) & (mul_34_17_n_10789 | mul_34_17_n_10464));
 assign mul_34_17_n_10806 = ((mul_34_17_n_10599 | mul_34_17_n_10534) & (mul_34_17_n_10790 | mul_34_17_n_10592));
 assign mul_34_17_n_10803 = ~(mul_34_17_n_10788 | mul_34_17_n_10854);
 assign mul_34_17_n_10802 = ~(mul_34_17_n_10789 | mul_34_17_n_10550);
 assign mul_34_17_n_10801 = ~(mul_34_17_n_10785 | mul_34_17_n_10722);
 assign mul_34_17_n_10805 = ~(mul_34_17_n_10789 | mul_34_17_n_10501);
 assign mul_34_17_n_10800 = ~(mul_34_17_n_10786 & mul_34_17_n_10704);
 assign mul_34_17_n_10799 = ((mul_34_17_n_10827 & mul_34_17_n_10284) | ((mul_34_17_n_10827 & mul_34_17_n_10893)
    | (mul_34_17_n_10893 & mul_34_17_n_10284)));
 assign mul_34_17_n_10798 = ~(mul_34_17_n_10787 & mul_34_17_n_10779);
 assign mul_34_17_n_10804 = ~(mul_34_17_n_10791 & mul_34_17_n_10783);
 assign asc001_58_ = ~(mul_34_17_n_10777 ^ mul_34_17_n_10447);
 assign mul_34_17_n_10797 = ((mul_34_17_n_10896 & mul_34_17_n_10897) | (mul_34_17_n_10784 & mul_34_17_n_10646));
 assign asc001_65_ = ~(mul_34_17_n_10778 ^ mul_34_17_n_10584);
 assign mul_34_17_n_10796 = ((mul_34_17_n_10440 | mul_34_17_n_10916) & (mul_34_17_n_10783 | mul_34_17_n_10610));
 assign mul_34_17_n_10795 = ~(mul_34_17_n_10383 | (mul_34_17_n_10340 | (mul_34_17_n_10550 | mul_34_17_n_10789)));
 assign mul_34_17_n_10794 = ((mul_34_17_n_10671 & mul_34_17_n_10306) | (mul_34_17_n_10776 & mul_34_17_n_10613));
 assign asc001_66_ = ~(mul_34_17_n_10284 ^ mul_34_17_n_10450);
 assign mul_34_17_n_10793 = ~(mul_34_17_n_10782 & (mul_34_17_n_10678 & (mul_34_17_n_10714 & mul_34_17_n_10395)));
 assign mul_34_17_n_10792 = ~(mul_34_17_n_10780 & (mul_34_17_n_10857 & (mul_34_17_n_10721 & mul_34_17_n_10459)));
 assign mul_34_17_n_10788 = ~(mul_34_17_n_10783 | mul_34_17_n_10647);
 assign mul_34_17_n_10787 = ~(mul_34_17_n_10776 & mul_34_17_n_10611);
 assign asc001_60_ = (mul_34_17_n_10371 ^ mul_34_17_n_10766);
 assign mul_34_17_n_10786 = ~(mul_34_17_n_10781 | mul_34_17_n_10293);
 assign mul_34_17_n_10785 = ((mul_34_17_n_10876 & mul_34_17_n_10775) | ((mul_34_17_n_10876 & mul_34_17_n_11017)
    | (mul_34_17_n_11017 & mul_34_17_n_10775)));
 assign mul_34_17_n_10791 = ~(mul_34_17_n_10750 & (mul_34_17_n_10645 & (mul_34_17_n_10676 & mul_34_17_n_10621)));
 assign mul_34_17_n_10790 = ~(mul_34_17_n_10784 | mul_34_17_n_10697);
 assign mul_34_17_n_10789 = ~(mul_34_17_n_10776 | mul_34_17_n_10732);
 assign asc001_52_ = ~(mul_34_17_n_10770 ^ mul_34_17_n_10332);
 assign asc001_56_ = ~(mul_34_17_n_10769 ^ mul_34_17_n_10324);
 assign asc001_54_ = ~(mul_34_17_n_10767 ^ mul_34_17_n_10325);
 assign asc001_53_ = ~(mul_34_17_n_10762 ^ mul_34_17_n_10491);
 assign asc001_57_ = ~(mul_34_17_n_10768 ^ mul_34_17_n_10547);
 assign asc001_51_ = ~(mul_34_17_n_10761 ^ mul_34_17_n_10444);
 assign asc001_50_ = ~(mul_34_17_n_10763 ^ mul_34_17_n_10416);
 assign asc001_49_ = ~(mul_34_17_n_10764 ^ mul_34_17_n_10452);
 assign mul_34_17_n_10782 = ~(mul_34_17_n_10771 & mul_34_17_n_10588);
 assign mul_34_17_n_10781 = ~(mul_34_17_n_10772 | mul_34_17_n_10303);
 assign mul_34_17_n_10780 = ~(mul_34_17_n_10760 & (mul_34_17_n_10588 & (mul_34_17_n_10357 & mul_34_17_n_11024)));
 assign mul_34_17_n_10779 = ~(mul_34_17_n_10765 | mul_34_17_n_10467);
 assign mul_34_17_n_10778 = ((mul_34_17_n_10593 & mul_34_17_n_10750) | ((mul_34_17_n_10593 & mul_34_17_n_10364)
    | (mul_34_17_n_10364 & mul_34_17_n_10750)));
 assign mul_34_17_n_10784 = ~(mul_34_17_n_10774 | mul_34_17_n_10644);
 assign mul_34_17_n_10777 = ~(mul_34_17_n_10775 | mul_34_17_n_10710);
 assign mul_34_17_n_10783 = ~(mul_34_17_n_10755 | (mul_34_17_n_10681 | (mul_34_17_n_10624 | mul_34_17_n_10517)));
 assign asc001_43_ = ~(mul_34_17_n_10745 ^ mul_34_17_n_10422);
 assign asc001_46_ = ~(mul_34_17_n_10754 ^ mul_34_17_n_10323);
 assign asc001_45_ = ~(mul_34_17_n_10743 ^ mul_34_17_n_10428);
 assign asc001_44_ = ~(mul_34_17_n_10752 ^ mul_34_17_n_10495);
 assign asc001_55_ = ~(mul_34_17_n_10744 ^ mul_34_17_n_10430);
 assign asc001_42_ = ~(mul_34_17_n_10753 ^ mul_34_17_n_10330);
 assign asc001_41_ = ~(mul_34_17_n_10746 ^ mul_34_17_n_10418);
 assign asc001_64_ = ~(mul_34_17_n_10750 ^ mul_34_17_n_10659);
 assign mul_34_17_n_10776 = ~(mul_34_17_n_10749 | (mul_34_17_n_10644 | (mul_34_17_n_10656 | mul_34_17_n_10632)));
 assign mul_34_17_n_10773 = ~(mul_34_17_n_10757 & mul_34_17_n_11041);
 assign mul_34_17_n_10772 = ~(mul_34_17_n_10751 | mul_34_17_n_10665);
 assign mul_34_17_n_10771 = ~(mul_34_17_n_10742 | (mul_34_17_n_10590 | (mul_34_17_n_10465 | mul_34_17_n_10339)));
 assign mul_34_17_n_10770 = ~(mul_34_17_n_10756 | mul_34_17_n_10641);
 assign mul_34_17_n_10775 = ~(mul_34_17_n_10742 | (mul_34_17_n_10590 | (mul_34_17_n_10510 | mul_34_17_n_11022)));
 assign mul_34_17_n_10769 = ~(mul_34_17_n_10760 | mul_34_17_n_10683);
 assign mul_34_17_n_10774 = ~(mul_34_17_n_10750 & mul_34_17_n_10657);
 assign mul_34_17_n_10768 = ~(mul_34_17_n_10700 | mul_34_17_n_10758);
 assign mul_34_17_n_10767 = ~(mul_34_17_n_10689 | mul_34_17_n_10747);
 assign mul_34_17_n_10766 = ~(mul_34_17_n_10751 | mul_34_17_n_10703);
 assign asc001_48_ = ~(mul_34_17_n_10742 ^ mul_34_17_n_10456);
 assign asc001_35_ = (mul_34_17_n_10929 ^ mul_34_17_n_10725);
 assign asc001_37_ = ~(mul_34_17_n_10727 ^ mul_34_17_n_10871);
 assign asc001_38_ = ~(mul_34_17_n_10733 ^ mul_34_17_n_10320);
 assign mul_34_17_n_10765 = ((mul_34_17_n_10671 & mul_34_17_n_10384) | (mul_34_17_n_10732 & mul_34_17_n_10611));
 assign asc001_39_ = (mul_34_17_n_11021 ^ mul_34_17_n_10734);
 assign asc001_47_ = ~(mul_34_17_n_10726 ^ mul_34_17_n_10493);
 assign mul_34_17_n_10764 = ((mul_34_17_n_10875 & mul_34_17_n_10741) | ((mul_34_17_n_10875 & mul_34_17_n_11019)
    | (mul_34_17_n_11019 & mul_34_17_n_10741)));
 assign mul_34_17_n_10763 = ((mul_34_17_n_10487 | mul_34_17_n_10342) & (mul_34_17_n_10742 | mul_34_17_n_10484));
 assign mul_34_17_n_10762 = ~(mul_34_17_n_10690 | mul_34_17_n_10759);
 assign mul_34_17_n_10761 = ~(mul_34_17_n_10691 | mul_34_17_n_10748);
 assign mul_34_17_n_10759 = ~(mul_34_17_n_10738 & mul_34_17_n_10843);
 assign mul_34_17_n_10758 = ~(mul_34_17_n_10740 & mul_34_17_n_10882);
 assign mul_34_17_n_10757 = ~(mul_34_17_n_10732 & mul_34_17_n_10613);
 assign mul_34_17_n_10756 = ~(mul_34_17_n_10742 | mul_34_17_n_10551);
 assign mul_34_17_n_10755 = ~(mul_34_17_n_10559 | (mul_34_17_n_10383 | (mul_34_17_n_10550 | mul_34_17_n_10731)));
 assign mul_34_17_n_10754 = ~(mul_34_17_n_10736 | mul_34_17_n_10653);
 assign mul_34_17_n_10753 = ~(mul_34_17_n_10739 | mul_34_17_n_10505);
 assign mul_34_17_n_10752 = ~(mul_34_17_n_10735 | mul_34_17_n_10609);
 assign mul_34_17_n_10760 = ~(mul_34_17_n_10742 | mul_34_17_n_10590);
 assign mul_34_17_n_10749 = ~mul_34_17_n_10750;
 assign asc001_40_ = ~(mul_34_17_n_10723 ^ mul_34_17_n_10417);
 assign mul_34_17_n_10748 = ~((mul_34_17_n_10859 | mul_34_17_n_10858) & (mul_34_17_n_10717 | mul_34_17_n_10539));
 assign mul_34_17_n_10747 = ~(mul_34_17_n_10737 & mul_34_17_n_10554);
 assign mul_34_17_n_10751 = ~(mul_34_17_n_10742 | mul_34_17_n_10625);
 assign mul_34_17_n_10746 = ((mul_34_17_n_10867 & mul_34_17_n_10723) | ((mul_34_17_n_10867 & mul_34_17_n_10860)
    | (mul_34_17_n_10860 & mul_34_17_n_10723)));
 assign mul_34_17_n_10745 = ~(mul_34_17_n_10713 & (mul_34_17_n_11035 & (mul_34_17_n_10639 & mul_34_17_n_10570)));
 assign mul_34_17_n_10744 = ~(mul_34_17_n_10685 & (mul_34_17_n_10883 & (mul_34_17_n_10670 & mul_34_17_n_10730)));
 assign mul_34_17_n_10743 = ~(mul_34_17_n_10728 & mul_34_17_n_10655);
 assign mul_34_17_n_10750 = ~(mul_34_17_n_10682 & (mul_34_17_n_10586 & (mul_34_17_n_10701 & mul_34_17_n_10729)));
 assign mul_34_17_n_10741 = ~mul_34_17_n_10742;
 assign mul_34_17_n_10740 = ~(mul_34_17_n_10718 & mul_34_17_n_10648);
 assign mul_34_17_n_10739 = ~(mul_34_17_n_10723 | mul_34_17_n_10469);
 assign mul_34_17_n_10738 = ~(mul_34_17_n_10718 & mul_34_17_n_10614);
 assign mul_34_17_n_10737 = ~(mul_34_17_n_10718 & mul_34_17_n_10615);
 assign mul_34_17_n_10736 = ~(mul_34_17_n_10716 & mul_34_17_n_10553);
 assign mul_34_17_n_10735 = ~(mul_34_17_n_10723 | mul_34_17_n_10504);
 assign mul_34_17_n_10734 = ~(mul_34_17_n_10724 | mul_34_17_n_10480);
 assign mul_34_17_n_10733 = ~(mul_34_17_n_10719 | mul_34_17_n_11248);
 assign mul_34_17_n_10742 = ~(mul_34_17_n_10680 | mul_34_17_n_10718);
 assign mul_34_17_n_10732 = ~mul_34_17_n_10731;
 assign mul_34_17_n_10730 = ~(mul_34_17_n_10718 & mul_34_17_n_10597);
 assign asc001_33_ = (mul_34_17_n_10869 ^ mul_34_17_n_10699);
 assign mul_34_17_n_10729 = ~(mul_34_17_n_10718 & mul_34_17_n_10658);
 assign asc001_34_ = ~(mul_34_17_n_10702 ^ mul_34_17_n_11028);
 assign mul_34_17_n_10728 = ((mul_34_17_n_10386 | mul_34_17_n_10379) & (mul_34_17_n_10706 | mul_34_17_n_10581));
 assign asc001_36_ = ~(mul_34_17_n_10709 ^ mul_34_17_n_10443);
 assign mul_34_17_n_10727 = ((mul_34_17_n_10928 & mul_34_17_n_10709) | ((mul_34_17_n_10928 & mul_34_17_n_10840)
    | (mul_34_17_n_10840 & mul_34_17_n_10709)));
 assign mul_34_17_n_10726 = ~(mul_34_17_n_10638 & (mul_34_17_n_10909 & (mul_34_17_n_10650 & mul_34_17_n_10715)));
 assign mul_34_17_n_10725 = ((mul_34_17_n_10834 | mul_34_17_n_10865) & (mul_34_17_n_10702 | mul_34_17_n_11044));
 assign mul_34_17_n_10731 = ~(mul_34_17_n_10705 | (mul_34_17_n_10476 | (mul_34_17_n_10654 | mul_34_17_n_10519)));
 assign mul_34_17_n_10724 = ~mul_34_17_n_10720;
 assign mul_34_17_n_10722 = ~(mul_34_17_n_10711 | mul_34_17_n_10378);
 assign mul_34_17_n_10721 = ~(mul_34_17_n_10703 & mul_34_17_n_10466);
 assign mul_34_17_n_10720 = ~(mul_34_17_n_10709 & mul_34_17_n_10407);
 assign mul_34_17_n_10719 = ~(mul_34_17_n_10708 | mul_34_17_n_10841);
 assign mul_34_17_n_10723 = ~(mul_34_17_n_10707 | mul_34_17_n_10607);
 assign mul_34_17_n_10717 = ~mul_34_17_n_10718;
 assign mul_34_17_n_10716 = ~(mul_34_17_n_10707 & mul_34_17_n_10580);
 assign mul_34_17_n_10715 = ~(mul_34_17_n_10707 & mul_34_17_n_10596);
 assign mul_34_17_n_10714 = ((mul_34_17_n_10513 | mul_34_17_n_10339) & (mul_34_17_n_10694 | mul_34_17_n_10530));
 assign mul_34_17_n_10713 = ~(mul_34_17_n_10707 & mul_34_17_n_10540);
 assign mul_34_17_n_10712 = ((mul_34_17_n_10619 & mul_34_17_n_10345) | (mul_34_17_n_10697 & mul_34_17_n_10646));
 assign mul_34_17_n_10718 = ~(mul_34_17_n_10688 | (mul_34_17_n_10489 | (mul_34_17_n_10485 | mul_34_17_n_10601)));
 assign mul_34_17_n_10711 = ~mul_34_17_n_10710;
 assign mul_34_17_n_10708 = ~mul_34_17_n_10709;
 assign mul_34_17_n_10706 = ~mul_34_17_n_10707;
 assign mul_34_17_n_10705 = ~(mul_34_17_n_10696 | mul_34_17_n_10632);
 assign mul_34_17_n_10704 = ~(mul_34_17_n_10695 & mul_34_17_n_11024);
 assign mul_34_17_n_10710 = ~(mul_34_17_n_10692 & mul_34_17_n_10594);
 assign mul_34_17_n_10709 = ~(mul_34_17_n_10698 & mul_34_17_n_10477);
 assign mul_34_17_n_10707 = ~(mul_34_17_n_10698 | mul_34_17_n_10485);
 assign mul_34_17_n_10701 = ~((mul_34_17_n_10683 & mul_34_17_n_10630) | (mul_34_17_n_10680 & mul_34_17_n_10658));
 assign mul_34_17_n_10700 = ((mul_34_17_n_10683 & mul_34_17_n_10291) | (mul_34_17_n_10680 & mul_34_17_n_10648));
 assign asc001_32_ = (mul_34_17_n_11029 ^ mul_34_17_n_10688);
 assign mul_34_17_n_10699 = ~((mul_34_17_n_10825 & mul_34_17_n_11036) | (mul_34_17_n_10687 & mul_34_17_n_11030));
 assign mul_34_17_n_10703 = ~(mul_34_17_n_10694 & mul_34_17_n_10666);
 assign mul_34_17_n_10702 = ~(mul_34_17_n_10693 | mul_34_17_n_10317);
 assign mul_34_17_n_10697 = ~mul_34_17_n_10696;
 assign mul_34_17_n_10695 = ~mul_34_17_n_10694;
 assign mul_34_17_n_10693 = ~(mul_34_17_n_10688 | mul_34_17_n_10402);
 assign mul_34_17_n_10692 = ~(mul_34_17_n_10683 & mul_34_17_n_10564);
 assign mul_34_17_n_10698 = ~(mul_34_17_n_10687 & mul_34_17_n_10488);
 assign mul_34_17_n_10696 = ~(mul_34_17_n_10686 | mul_34_17_n_10651);
 assign mul_34_17_n_10694 = ~(mul_34_17_n_10683 & mul_34_17_n_10588);
 assign mul_34_17_n_10691 = ~((mul_34_17_n_10506 | mul_34_17_n_10346) & (mul_34_17_n_10679 | mul_34_17_n_10539));
 assign mul_34_17_n_10690 = ((mul_34_17_n_10641 & mul_34_17_n_10304) | (mul_34_17_n_10680 & mul_34_17_n_10614));
 assign mul_34_17_n_10689 = ((mul_34_17_n_10641 & mul_34_17_n_10526) | (mul_34_17_n_10680 & mul_34_17_n_10615));
 assign asc001_30_ = ~(mul_34_17_n_10674 ^ mul_34_17_n_10333);
 assign asc001_29_ = ~(mul_34_17_n_10675 ^ mul_34_17_n_10968);
 assign mul_34_17_n_10687 = ~mul_34_17_n_10688;
 assign mul_34_17_n_10686 = ~(mul_34_17_n_10673 | mul_34_17_n_10644);
 assign mul_34_17_n_10685 = ~(mul_34_17_n_10680 & mul_34_17_n_10597);
 assign mul_34_17_n_10684 = ~(mul_34_17_n_10672 | mul_34_17_n_10454);
 assign mul_34_17_n_10688 = ~(mul_34_17_n_10652 | mul_34_17_n_10677);
 assign mul_34_17_n_10682 = ~((mul_34_17_n_10847 & mul_34_17_n_10886) | (mul_34_17_n_10665 & mul_34_17_n_10512));
 assign mul_34_17_n_10681 = ~(mul_34_17_n_10672 | mul_34_17_n_10612);
 assign asc001_31_ = ~(mul_34_17_n_10649 ^ mul_34_17_n_10992);
 assign mul_34_17_n_10683 = ~(mul_34_17_n_10669 & mul_34_17_n_10626);
 assign mul_34_17_n_10679 = ~mul_34_17_n_10680;
 assign mul_34_17_n_10678 = ~(mul_34_17_n_10665 & mul_34_17_n_10529);
 assign mul_34_17_n_10677 = ~(mul_34_17_n_10663 & mul_34_17_n_10991);
 assign mul_34_17_n_10676 = ~(mul_34_17_n_10656 | mul_34_17_n_10632);
 assign mul_34_17_n_10675 = ~(mul_34_17_n_10668 & mul_34_17_n_10969);
 assign mul_34_17_n_10674 = ~(mul_34_17_n_10660 & mul_34_17_n_11251);
 assign mul_34_17_n_10680 = ~(mul_34_17_n_10627 & (mul_34_17_n_10549 & (mul_34_17_n_10637 & mul_34_17_n_10604)));
 assign mul_34_17_n_10671 = ~mul_34_17_n_10672;
 assign mul_34_17_n_10670 = ((mul_34_17_n_10554 | mul_34_17_n_10881) & (mul_34_17_n_10640 | mul_34_17_n_10582));
 assign mul_34_17_n_10669 = ((mul_34_17_n_11043 | mul_34_17_n_11008) & (mul_34_17_n_10640 | mul_34_17_n_10557));
 assign asc001_27_ = (mul_34_17_n_10846 ^ mul_34_17_n_10634);
 assign asc001_28_ = ~(mul_34_17_n_10642 ^ mul_34_17_n_10327);
 assign mul_34_17_n_10673 = ~(mul_34_17_n_10664 | mul_34_17_n_10565);
 assign mul_34_17_n_10672 = ~(mul_34_17_n_10662 | mul_34_17_n_10321);
 assign mul_34_17_n_10668 = ~mul_34_17_n_10661;
 assign mul_34_17_n_10666 = ~mul_34_17_n_10665;
 assign mul_34_17_n_10664 = ~(mul_34_17_n_10633 | mul_34_17_n_10563);
 assign mul_34_17_n_10663 = ~(mul_34_17_n_10628 & mul_34_17_n_10308);
 assign mul_34_17_n_10662 = ~(mul_34_17_n_10631 | mul_34_17_n_10358);
 assign mul_34_17_n_10661 = ~(mul_34_17_n_10642 | mul_34_17_n_10967);
 assign mul_34_17_n_10660 = ~(mul_34_17_n_10643 & mul_34_17_n_10403);
 assign mul_34_17_n_10667 = ~(mul_34_17_n_10623 | mul_34_17_n_10605);
 assign mul_34_17_n_10659 = ~(mul_34_17_n_10593 ^ mul_34_17_n_10364);
 assign mul_34_17_n_10665 = ~(mul_34_17_n_10636 & mul_34_17_n_10548);
 assign mul_34_17_n_10657 = ~mul_34_17_n_10656;
 assign mul_34_17_n_10655 = ((mul_34_17_n_10608 | mul_34_17_n_10472) & (mul_34_17_n_10606 | mul_34_17_n_10581));
 assign mul_34_17_n_10654 = ~(mul_34_17_n_10599 | (mul_34_17_n_10534 | (mul_34_17_n_10470 | mul_34_17_n_10344)));
 assign mul_34_17_n_10653 = ((mul_34_17_n_10609 & mul_34_17_n_10524) | (mul_34_17_n_10580 & mul_34_17_n_10607));
 assign mul_34_17_n_10652 = ~((mul_34_17_n_10478 | mul_34_17_n_10993) & (mul_34_17_n_10616 | mul_34_17_n_10993));
 assign mul_34_17_n_10651 = ((mul_34_17_n_10556 & mul_34_17_n_10368) | ((mul_34_17_n_10556 & mul_34_17_n_10538)
    | (mul_34_17_n_10538 & mul_34_17_n_10368)));
 assign mul_34_17_n_10650 = ((mul_34_17_n_10553 | mul_34_17_n_10908) & (mul_34_17_n_10608 | mul_34_17_n_10583));
 assign mul_34_17_n_10649 = ~(mul_34_17_n_10635 | mul_34_17_n_10628);
 assign mul_34_17_n_10658 = ~(mul_34_17_n_10629 | mul_34_17_n_10590);
 assign mul_34_17_n_10656 = ~((mul_34_17_n_10509 | mul_34_17_n_10399) & (mul_34_17_n_10593 | mul_34_17_n_10364));
 assign mul_34_17_n_10645 = ~mul_34_17_n_10644;
 assign mul_34_17_n_10643 = ~mul_34_17_n_10642;
 assign mul_34_17_n_10640 = ~mul_34_17_n_10641;
 assign mul_34_17_n_10639 = ~(mul_34_17_n_10607 & mul_34_17_n_10540);
 assign mul_34_17_n_10638 = ~(mul_34_17_n_10596 & mul_34_17_n_10607);
 assign mul_34_17_n_10637 = ~(mul_34_17_n_10609 & mul_34_17_n_10579);
 assign mul_34_17_n_10636 = ~(mul_34_17_n_10595 & mul_34_17_n_10515);
 assign mul_34_17_n_10635 = ~(mul_34_17_n_10616 & mul_34_17_n_10478);
 assign mul_34_17_n_10634 = ~(mul_34_17_n_10602 | mul_34_17_n_10935);
 assign mul_34_17_n_10648 = ~(mul_34_17_n_10590 | mul_34_17_n_11022);
 assign mul_34_17_n_10647 = ~(mul_34_17_n_10598 & mul_34_17_n_10313);
 assign mul_34_17_n_10646 = ~(mul_34_17_n_10592 | mul_34_17_n_10344);
 assign mul_34_17_n_10633 = ~(mul_34_17_n_10593 & mul_34_17_n_10364);
 assign mul_34_17_n_10644 = ~(mul_34_17_n_10600 & mul_34_17_n_10367);
 assign mul_34_17_n_10642 = ~(mul_34_17_n_10618 | mul_34_17_n_10560);
 assign mul_34_17_n_10641 = ~(mul_34_17_n_10587 & mul_34_17_n_10462);
 assign mul_34_17_n_10632 = ~mul_34_17_n_10622;
 assign mul_34_17_n_10630 = ~mul_34_17_n_10629;
 assign mul_34_17_n_10627 = ~(mul_34_17_n_10541 & (mul_34_17_n_10524 & (mul_34_17_n_10503 & mul_34_17_n_10607)));
 assign asc001_26_ = ~(mul_34_17_n_10567 ^ mul_34_17_n_10936);
 assign mul_34_17_n_10626 = ((mul_34_17_n_10883 | mul_34_17_n_10839) & (mul_34_17_n_10554 | mul_34_17_n_10410));
 assign mul_34_17_n_10625 = ~(mul_34_17_n_10589 & mul_34_17_n_10588);
 assign mul_34_17_n_10624 = ((mul_34_17_n_10536 & mul_34_17_n_10353) | (mul_34_17_n_10558 & mul_34_17_n_10467));
 assign mul_34_17_n_10623 = ~(mul_34_17_n_10591 | mul_34_17_n_10578);
 assign mul_34_17_n_10622 = ~(mul_34_17_n_10577 | (mul_34_17_n_10534 | (mul_34_17_n_10470 | mul_34_17_n_10344)));
 assign mul_34_17_n_10631 = ~(mul_34_17_n_10603 | mul_34_17_n_10398);
 assign mul_34_17_n_10629 = ~(mul_34_17_n_10588 & mul_34_17_n_10512);
 assign mul_34_17_n_10621 = ~(mul_34_17_n_10612 | mul_34_17_n_10550);
 assign mul_34_17_n_10628 = ~(mul_34_17_n_10617 | mul_34_17_n_10481);
 assign mul_34_17_n_10620 = (mul_34_17_n_10556 ^ mul_34_17_n_10538);
 assign mul_34_17_n_10619 = ~(mul_34_17_n_10599 | mul_34_17_n_10534);
 assign mul_34_17_n_10618 = ~mul_34_17_n_10617;
 assign mul_34_17_n_10608 = ~mul_34_17_n_10609;
 assign mul_34_17_n_10606 = ~mul_34_17_n_10607;
 assign mul_34_17_n_10605 = ~(mul_34_17_n_10568 & mul_34_17_n_10408);
 assign mul_34_17_n_10604 = ~(mul_34_17_n_10552 & mul_34_17_n_10541);
 assign mul_34_17_n_10603 = ~(mul_34_17_n_10561 | mul_34_17_n_10381);
 assign mul_34_17_n_10602 = ~(mul_34_17_n_10573 | mul_34_17_n_10319);
 assign mul_34_17_n_10617 = ~(mul_34_17_n_10569 | mul_34_17_n_10301);
 assign mul_34_17_n_10616 = ~(mul_34_17_n_10560 & mul_34_17_n_10482);
 assign mul_34_17_n_10615 = ~(mul_34_17_n_10551 | mul_34_17_n_10525);
 assign mul_34_17_n_10614 = ~(mul_34_17_n_10551 | mul_34_17_n_11038);
 assign mul_34_17_n_10613 = ~(mul_34_17_n_10550 | mul_34_17_n_10942);
 assign mul_34_17_n_10601 = ~(mul_34_17_n_10579 & mul_34_17_n_10503);
 assign mul_34_17_n_10612 = ~(mul_34_17_n_10558 & mul_34_17_n_10384);
 assign mul_34_17_n_10611 = ~(mul_34_17_n_10550 | mul_34_17_n_10383);
 assign mul_34_17_n_10610 = ~(mul_34_17_n_10575 & mul_34_17_n_10527);
 assign mul_34_17_n_10600 = ~(mul_34_17_n_10555 & mul_34_17_n_10537);
 assign mul_34_17_n_10609 = ~(mul_34_17_n_10571 & mul_34_17_n_10499);
 assign mul_34_17_n_10607 = ~(mul_34_17_n_10572 & mul_34_17_n_10521);
 assign mul_34_17_n_10595 = ~mul_34_17_n_10594;
 assign mul_34_17_n_10590 = ~mul_34_17_n_10589;
 assign mul_34_17_n_10599 = ~(mul_34_17_n_10543 | mul_34_17_n_10282);
 assign asc001_25_ = ~(mul_34_17_n_10516 ^ mul_34_17_n_10429);
 assign asc001_19_ = (mul_34_17_n_10961 ^ mul_34_17_n_10492);
 assign mul_34_17_n_10587 = ((mul_34_17_n_11007 | mul_34_17_n_10842) & (mul_34_17_n_10506 | mul_34_17_n_10420));
 assign mul_34_17_n_10586 = ((mul_34_17_n_10388 | mul_34_17_n_10395) & (mul_34_17_n_10513 | mul_34_17_n_10441));
 assign mul_34_17_n_10598 = ~(mul_34_17_n_10574 | mul_34_17_n_10578);
 assign mul_34_17_n_10597 = ~(mul_34_17_n_10551 | mul_34_17_n_10582);
 assign mul_34_17_n_10596 = ~(mul_34_17_n_10583 | mul_34_17_n_10504);
 assign mul_34_17_n_10594 = ((mul_34_17_n_10463 & mul_34_17_n_10392) | ((mul_34_17_n_10463 & mul_34_17_n_10882)
    | (mul_34_17_n_10882 & mul_34_17_n_10392)));
 assign mul_34_17_n_10593 = ~(mul_34_17_n_10494 ^ mul_34_17_n_11006);
 assign mul_34_17_n_10585 = ~(mul_34_17_n_10511 ^ mul_34_17_n_10436);
 assign mul_34_17_n_10584 = ~(mul_34_17_n_10509 ^ mul_34_17_n_10399);
 assign mul_34_17_n_10592 = ~(mul_34_17_n_10576 & mul_34_17_n_10533);
 assign mul_34_17_n_10591 = ~((mul_34_17_n_10913 & mul_34_17_n_10915) | (mul_34_17_n_10514 & mul_34_17_n_10302));
 assign mul_34_17_n_10589 = ~(mul_34_17_n_10557 | mul_34_17_n_10551);
 assign mul_34_17_n_10588 = ~(mul_34_17_n_10510 | (mul_34_17_n_11022 | (mul_34_17_n_10471 | mul_34_17_n_10378)));
 assign mul_34_17_n_10577 = ~mul_34_17_n_10576;
 assign mul_34_17_n_10575 = ~mul_34_17_n_10574;
 assign mul_34_17_n_10573 = ~(mul_34_17_n_10508 | mul_34_17_n_10522);
 assign mul_34_17_n_10572 = ~(mul_34_17_n_10518 | mul_34_17_n_10863);
 assign mul_34_17_n_10571 = ~(mul_34_17_n_10505 & mul_34_17_n_10460);
 assign mul_34_17_n_10570 = ~(mul_34_17_n_10505 & mul_34_17_n_10305);
 assign mul_34_17_n_10569 = ~(mul_34_17_n_10507 | mul_34_17_n_11005);
 assign mul_34_17_n_10568 = ~(mul_34_17_n_10531 & mul_34_17_n_10351);
 assign mul_34_17_n_10583 = ~(mul_34_17_n_10524 & mul_34_17_n_10288);
 assign mul_34_17_n_10567 = ~(mul_34_17_n_10507 & mul_34_17_n_10520);
 assign mul_34_17_n_10582 = ~(mul_34_17_n_10526 & mul_34_17_n_10290);
 assign mul_34_17_n_10581 = ~(mul_34_17_n_10503 & mul_34_17_n_10473);
 assign mul_34_17_n_10580 = ~(mul_34_17_n_10504 | mul_34_17_n_10523);
 assign mul_34_17_n_10579 = ~(mul_34_17_n_10475 | (mul_34_17_n_10908 | (mul_34_17_n_10472 | mul_34_17_n_10905)));
 assign mul_34_17_n_10566 = ~(mul_34_17_n_10534 | mul_34_17_n_10282);
 assign mul_34_17_n_10565 = ~((mul_34_17_n_11004 & mul_34_17_n_11050) | (mul_34_17_n_10490 & mul_34_17_n_10412));
 assign mul_34_17_n_10578 = ~(mul_34_17_n_10527 & mul_34_17_n_10351);
 assign mul_34_17_n_10564 = ~(mul_34_17_n_10510 | mul_34_17_n_11022);
 assign mul_34_17_n_10576 = ~(mul_34_17_n_10511 & mul_34_17_n_10436);
 assign mul_34_17_n_10563 = ~(mul_34_17_n_10509 | mul_34_17_n_10399);
 assign mul_34_17_n_10574 = ~((mul_34_17_n_10913 | mul_34_17_n_10915) & (mul_34_17_n_10435 | mul_34_17_n_10362));
 assign mul_34_17_n_10562 = ~mul_34_17_n_10561;
 assign mul_34_17_n_10559 = ~mul_34_17_n_10558;
 assign mul_34_17_n_10556 = ~mul_34_17_n_10555;
 assign mul_34_17_n_10553 = ~mul_34_17_n_10552;
 assign mul_34_17_n_10550 = ~mul_34_17_n_10542;
 assign mul_34_17_n_10549 = ((mul_34_17_n_10382 & mul_34_17_n_10359) | ((mul_34_17_n_10382 & mul_34_17_n_10909)
    | (mul_34_17_n_10909 & mul_34_17_n_10359)));
 assign mul_34_17_n_10548 = ((mul_34_17_n_10411 | mul_34_17_n_10406) & (mul_34_17_n_10471 | mul_34_17_n_10355));
 assign asc001_18_ = ~(mul_34_17_n_10426 ^ mul_34_17_n_10396);
 assign asc001_21_ = ~(mul_34_17_n_10423 ^ mul_34_17_n_10956);
 assign asc001_22_ = ~(mul_34_17_n_10458 ^ mul_34_17_n_10965);
 assign asc001_24_ = ~(mul_34_17_n_10419 ^ mul_34_17_n_10376);
 assign mul_34_17_n_10561 = ~((mul_34_17_n_10925 & mul_34_17_n_10950) | (mul_34_17_n_10474 & mul_34_17_n_10298));
 assign mul_34_17_n_10560 = ~(mul_34_17_n_10394 | (mul_34_17_n_11014 | (mul_34_17_n_11005 | mul_34_17_n_10377)));
 assign mul_34_17_n_10547 = ~(mul_34_17_n_10510 | mul_34_17_n_10502);
 assign mul_34_17_n_10558 = ~(mul_34_17_n_10535 | mul_34_17_n_10340);
 assign mul_34_17_n_10546 = ~(mul_34_17_n_10532 & mul_34_17_n_10527);
 assign mul_34_17_n_10557 = ~(mul_34_17_n_10526 & mul_34_17_n_10409);
 assign mul_34_17_n_10545 = (mul_34_17_n_10435 ^ mul_34_17_n_10363);
 assign mul_34_17_n_10555 = ~(mul_34_17_n_10427 ^ mul_34_17_n_10890);
 assign mul_34_17_n_10544 = ~(mul_34_17_n_10953 ^ mul_34_17_n_10438);
 assign mul_34_17_n_10554 = ((mul_34_17_n_10385 & mul_34_17_n_10360) | ((mul_34_17_n_10385 & mul_34_17_n_10843)
    | (mul_34_17_n_10843 & mul_34_17_n_10360)));
 assign mul_34_17_n_10552 = ~((mul_34_17_n_10945 | mul_34_17_n_10906) & (mul_34_17_n_10421 | mul_34_17_n_10905));
 assign mul_34_17_n_10543 = ~(mul_34_17_n_10511 | mul_34_17_n_10436);
 assign mul_34_17_n_10551 = ~(mul_34_17_n_10361 & (mul_34_17_n_10347 & (mul_34_17_n_10343 & mul_34_17_n_10874)));
 assign mul_34_17_n_10542 = ~(mul_34_17_n_10464 | (mul_34_17_n_10994 | (mul_34_17_n_10358 | mul_34_17_n_10381)));
 assign mul_34_17_n_10537 = ~mul_34_17_n_10538;
 assign mul_34_17_n_10536 = ~mul_34_17_n_10535;
 assign mul_34_17_n_10533 = ~mul_34_17_n_10534;
 assign mul_34_17_n_10532 = ~mul_34_17_n_10531;
 assign mul_34_17_n_10530 = ~mul_34_17_n_10529;
 assign mul_34_17_n_10528 = ~mul_34_17_n_10527;
 assign mul_34_17_n_10525 = ~mul_34_17_n_10526;
 assign mul_34_17_n_10523 = ~mul_34_17_n_10524;
 assign mul_34_17_n_10522 = ~(mul_34_17_n_10479 | mul_34_17_n_11014);
 assign mul_34_17_n_10521 = ~(mul_34_17_n_10480 & mul_34_17_n_10315);
 assign mul_34_17_n_10520 = ~(mul_34_17_n_10457 & mul_34_17_n_10376);
 assign mul_34_17_n_10519 = ~(mul_34_17_n_10470 | mul_34_17_n_10349);
 assign mul_34_17_n_10518 = ~(mul_34_17_n_10485 | mul_34_17_n_10477);
 assign mul_34_17_n_10517 = ~(mul_34_17_n_10439 | mul_34_17_n_10953);
 assign mul_34_17_n_10516 = ~(mul_34_17_n_10479 & mul_34_17_n_10352);
 assign mul_34_17_n_10541 = ~(mul_34_17_n_10475 | mul_34_17_n_10908);
 assign mul_34_17_n_10540 = ~(mul_34_17_n_10469 | mul_34_17_n_10872);
 assign mul_34_17_n_10539 = ~(mul_34_17_n_10483 & mul_34_17_n_10347);
 assign mul_34_17_n_10515 = ~(mul_34_17_n_10471 | mul_34_17_n_10378);
 assign mul_34_17_n_10538 = ~(mul_34_17_n_10433 & mul_34_17_n_10894);
 assign mul_34_17_n_10535 = ~(mul_34_17_n_10438 | mul_34_17_n_10297);
 assign mul_34_17_n_10514 = ~(mul_34_17_n_10434 | mul_34_17_n_10363);
 assign mul_34_17_n_10534 = ~(mul_34_17_n_10437 | mul_34_17_n_10365);
 assign mul_34_17_n_10531 = ~(mul_34_17_n_10440 | mul_34_17_n_10916);
 assign mul_34_17_n_10529 = ~(mul_34_17_n_10465 | mul_34_17_n_10339);
 assign mul_34_17_n_10527 = ~(mul_34_17_n_10440 & mul_34_17_n_10916);
 assign mul_34_17_n_10526 = ~(mul_34_17_n_10446 | mul_34_17_n_11038);
 assign mul_34_17_n_10524 = ~(mul_34_17_n_10472 | mul_34_17_n_10905);
 assign mul_34_17_n_10508 = ~mul_34_17_n_10507;
 assign mul_34_17_n_10503 = ~mul_34_17_n_10504;
 assign mul_34_17_n_10502 = ~(mul_34_17_n_10463 | mul_34_17_n_10392);
 assign mul_34_17_n_10501 = ~((mul_34_17_n_10925 | mul_34_17_n_10950) & (mul_34_17_n_10401 | mul_34_17_n_10405));
 assign mul_34_17_n_10500 = ~(mul_34_17_n_10468 | mul_34_17_n_10340);
 assign mul_34_17_n_10499 = ((mul_34_17_n_10939 & mul_34_17_n_11035) | ((mul_34_17_n_10939 & mul_34_17_n_10931)
    | (mul_34_17_n_10931 & mul_34_17_n_11035)));
 assign asc001_23_ = ~(mul_34_17_n_10322 ^ mul_34_17_n_10963);
 assign mul_34_17_n_10498 = ~(mul_34_17_n_10464 | mul_34_17_n_10474);
 assign mul_34_17_n_10497 = ~(mul_34_17_n_10470 | mul_34_17_n_10476);
 assign mul_34_17_n_10496 = ~(mul_34_17_n_10471 | mul_34_17_n_10424);
 assign mul_34_17_n_10495 = (mul_34_17_n_10379 ^ mul_34_17_n_10386);
 assign mul_34_17_n_10513 = ((mul_34_17_n_10885 & mul_34_17_n_10831) | ((mul_34_17_n_10885 & mul_34_17_n_10856)
    | (mul_34_17_n_10856 & mul_34_17_n_10831)));
 assign mul_34_17_n_10494 = ~(mul_34_17_n_10387 ^ mul_34_17_n_11000);
 assign mul_34_17_n_10512 = ~(mul_34_17_n_10441 | mul_34_17_n_10465);
 assign mul_34_17_n_10511 = ((mul_34_17_n_10289 & mul_34_17_n_10311) | ((mul_34_17_n_10289 & mul_34_17_n_11253)
    | (mul_34_17_n_11253 & mul_34_17_n_10311)));
 assign mul_34_17_n_10493 = ~(mul_34_17_n_10359 ^ mul_34_17_n_10382);
 assign mul_34_17_n_10510 = ~(mul_34_17_n_10413 | (mul_34_17_n_11049 | (mul_34_17_n_10880 | mul_34_17_n_10878)));
 assign mul_34_17_n_10492 = ((mul_34_17_n_10981 | mul_34_17_n_11015) & (mul_34_17_n_10396 | mul_34_17_n_10932));
 assign mul_34_17_n_10491 = (mul_34_17_n_10360 ^ mul_34_17_n_10385);
 assign mul_34_17_n_10509 = ~(mul_34_17_n_10490 & mul_34_17_n_10412);
 assign mul_34_17_n_10507 = ((mul_34_17_n_10937 | mul_34_17_n_10938) & (mul_34_17_n_10352 | mul_34_17_n_11014));
 assign mul_34_17_n_10506 = ~(mul_34_17_n_10486 & mul_34_17_n_10343);
 assign mul_34_17_n_10505 = ((mul_34_17_n_10861 & mul_34_17_n_10870) | (mul_34_17_n_10370 & mul_34_17_n_10862));
 assign mul_34_17_n_10504 = ~(mul_34_17_n_10390 & (mul_34_17_n_10305 & (mul_34_17_n_10397 & mul_34_17_n_10862)));
 assign mul_34_17_n_10489 = ~mul_34_17_n_10488;
 assign mul_34_17_n_10487 = ~mul_34_17_n_10486;
 assign mul_34_17_n_10484 = ~mul_34_17_n_10483;
 assign mul_34_17_n_10482 = ~mul_34_17_n_10481;
 assign mul_34_17_n_10473 = ~mul_34_17_n_10472;
 assign mul_34_17_n_10468 = ~mul_34_17_n_10467;
 assign mul_34_17_n_10466 = ~mul_34_17_n_10465;
 assign mul_34_17_n_10490 = ~(mul_34_17_n_10415 & mul_34_17_n_10387);
 assign mul_34_17_n_10488 = ~(mul_34_17_n_10402 | mul_34_17_n_10930);
 assign mul_34_17_n_10486 = ~(mul_34_17_n_10366 & mul_34_17_n_10873);
 assign mul_34_17_n_10462 = ~(mul_34_17_n_10348 & mul_34_17_n_10361);
 assign mul_34_17_n_10461 = ~(mul_34_17_n_10398 | mul_34_17_n_10381);
 assign mul_34_17_n_10460 = ~(mul_34_17_n_10391 | mul_34_17_n_10872);
 assign mul_34_17_n_10485 = ~(mul_34_17_n_10407 & mul_34_17_n_10315);
 assign mul_34_17_n_10483 = ~(mul_34_17_n_10369 | mul_34_17_n_10342);
 assign mul_34_17_n_10481 = ~(mul_34_17_n_10403 & mul_34_17_n_10294);
 assign mul_34_17_n_10480 = ~(mul_34_17_n_10335 & mul_34_17_n_11034);
 assign mul_34_17_n_10479 = ~(mul_34_17_n_10393 & mul_34_17_n_10376);
 assign mul_34_17_n_10478 = ~(mul_34_17_n_10373 | mul_34_17_n_10314);
 assign mul_34_17_n_10459 = ~(mul_34_17_n_10357 & mul_34_17_n_10293);
 assign mul_34_17_n_10477 = ~(mul_34_17_n_10336 | mul_34_17_n_10835);
 assign mul_34_17_n_10458 = ~(mul_34_17_n_10337 | mul_34_17_n_10957);
 assign mul_34_17_n_10457 = ~(mul_34_17_n_10394 | mul_34_17_n_11014);
 assign mul_34_17_n_10456 = (mul_34_17_n_10875 ^ mul_34_17_n_11019);
 assign mul_34_17_n_10455 = (mul_34_17_n_10941 ^ mul_34_17_n_10940);
 assign mul_34_17_n_10454 = ~(mul_34_17_n_10384 & mul_34_17_n_10341);
 assign mul_34_17_n_10476 = ~(mul_34_17_n_10331 | mul_34_17_n_10326);
 assign mul_34_17_n_10453 = (mul_34_17_n_10925 ^ mul_34_17_n_10950);
 assign mul_34_17_n_10452 = ~(mul_34_17_n_10366 & mul_34_17_n_10343);
 assign mul_34_17_n_10451 = ~(mul_34_17_n_10344 | mul_34_17_n_10350);
 assign mul_34_17_n_10450 = (mul_34_17_n_10827 ^ mul_34_17_n_10893);
 assign mul_34_17_n_10475 = ~(mul_34_17_n_10907 | (mul_34_17_n_11018 | (mul_34_17_n_10997 | mul_34_17_n_10828)));
 assign mul_34_17_n_10449 = ~(mul_34_17_n_10847 ^ mul_34_17_n_10886);
 assign mul_34_17_n_10448 = ~(mul_34_17_n_10338 & mul_34_17_n_10395);
 assign mul_34_17_n_10447 = ~(mul_34_17_n_10378 | mul_34_17_n_10356);
 assign mul_34_17_n_10446 = ~(mul_34_17_n_10850 | (mul_34_17_n_11002 | (mul_34_17_n_11023 | mul_34_17_n_10879)));
 assign mul_34_17_n_10445 = ~(mul_34_17_n_10408 & mul_34_17_n_10351);
 assign mul_34_17_n_10444 = (mul_34_17_n_11007 ^ mul_34_17_n_10842);
 assign mul_34_17_n_10443 = ~(mul_34_17_n_10928 ^ mul_34_17_n_10840);
 assign mul_34_17_n_10442 = ~(mul_34_17_n_10357 & mul_34_17_n_10857);
 assign mul_34_17_n_10474 = ~(mul_34_17_n_10400 | mul_34_17_n_10404);
 assign mul_34_17_n_10472 = ~(mul_34_17_n_10902 | (mul_34_17_n_10901 | (mul_34_17_n_10904 | mul_34_17_n_10900)));
 assign mul_34_17_n_10471 = ~(mul_34_17_n_10877 | (mul_34_17_n_10903 | (mul_34_17_n_11016 | mul_34_17_n_10832)));
 assign mul_34_17_n_10470 = ~(mul_34_17_n_10999 | (mul_34_17_n_11020 | (mul_34_17_n_10923 | mul_34_17_n_11031)));
 assign mul_34_17_n_10469 = ~(mul_34_17_n_10397 & mul_34_17_n_10862);
 assign mul_34_17_n_10467 = ~(mul_34_17_n_10414 & mul_34_17_n_10912);
 assign mul_34_17_n_10465 = ~(mul_34_17_n_10357 & mul_34_17_n_11024);
 assign mul_34_17_n_10464 = ~(mul_34_17_n_10401 | mul_34_17_n_10405);
 assign mul_34_17_n_10463 = ~(mul_34_17_n_10413 | mul_34_17_n_11049);
 assign mul_34_17_n_10439 = ~mul_34_17_n_10438;
 assign mul_34_17_n_10434 = ~mul_34_17_n_10435;
 assign asc001_14_ = ~(mul_34_17_n_10980 ^ mul_34_17_n_10989);
 assign asc001_11_ = ~(mul_34_17_n_10979 ^ mul_34_17_n_10852);
 assign asc001_8_ = ~(mul_34_17_n_10985 ^ mul_34_17_n_10976);
 assign asc001_7_ = ~(mul_34_17_n_11012 ^ mul_34_17_n_10975);
 assign asc001_5_ = ~(mul_34_17_n_11026 ^ mul_34_17_n_10987);
 assign asc001_6_ = ~(mul_34_17_n_10974 ^ mul_34_17_n_10986);
 assign asc001_4_ = ~(mul_34_17_n_11027 ^ mul_34_17_n_11039);
 assign asc001_3_ = ~(mul_34_17_n_11040 ^ mul_34_17_n_11048);
 assign asc001_1_ = ~(mul_34_17_n_10988 ^ mul_34_17_n_10943);
 assign asc001_12_ = ~(mul_34_17_n_11009 ^ mul_34_17_n_10982);
 assign mul_34_17_n_10433 = ((mul_34_17_n_10855 & mul_34_17_n_10889) | (mul_34_17_n_10891 & mul_34_17_n_10892));
 assign asc001_20_ = ~(mul_34_17_n_10960 ^ mul_34_17_n_11042);
 assign asc001_10_ = ~(mul_34_17_n_10977 ^ mul_34_17_n_10851);
 assign asc001_17_ = ~(mul_34_17_n_10927 ^ mul_34_17_n_10934);
 assign asc001_2_ = ~(mul_34_17_n_11037 ^ mul_34_17_n_11013);
 assign asc001_9_ = ~(mul_34_17_n_11010 ^ mul_34_17_n_10978);
 assign asc001_16_ = ~(mul_34_17_n_10837 ^ mul_34_17_n_10833);
 assign asc001_15_ = ~(mul_34_17_n_10973 ^ mul_34_17_n_10990);
 assign asc001_13_ = ~(mul_34_17_n_10984 ^ mul_34_17_n_11045);
 assign mul_34_17_n_10432 = ~(mul_34_17_n_10913 ^ mul_34_17_n_10915);
 assign mul_34_17_n_10441 = ~(mul_34_17_n_10389 & mul_34_17_n_10338);
 assign mul_34_17_n_10431 = ~(mul_34_17_n_10354 & mul_34_17_n_10341);
 assign mul_34_17_n_10430 = ~(mul_34_17_n_11043 ^ mul_34_17_n_11008);
 assign mul_34_17_n_10440 = ~(mul_34_17_n_10919 ^ mul_34_17_n_10917);
 assign mul_34_17_n_10429 = ~(mul_34_17_n_10937 ^ mul_34_17_n_10938);
 assign mul_34_17_n_10428 = ~(mul_34_17_n_10945 ^ mul_34_17_n_10906);
 assign mul_34_17_n_10427 = ~(mul_34_17_n_11253 ^ mul_34_17_n_11252);
 assign mul_34_17_n_10438 = (mul_34_17_n_10910 ^ mul_34_17_n_10954);
 assign mul_34_17_n_10426 = (mul_34_17_n_10981 ^ mul_34_17_n_11015);
 assign mul_34_17_n_10437 = ~(mul_34_17_n_10895 ^ mul_34_17_n_10898);
 assign mul_34_17_n_10436 = ~(mul_34_17_n_11033 ^ mul_34_17_n_10921);
 assign mul_34_17_n_10425 = ~(mul_34_17_n_11001 ^ mul_34_17_n_10920);
 assign mul_34_17_n_10424 = ~(mul_34_17_n_10411 | mul_34_17_n_10406);
 assign mul_34_17_n_10423 = ((mul_34_17_n_10962 & mul_34_17_n_10958) | (mul_34_17_n_10959 & mul_34_17_n_11042));
 assign mul_34_17_n_10435 = ~(mul_34_17_n_11032 ^ mul_34_17_n_10996);
 assign mul_34_17_n_10422 = ~(mul_34_17_n_10939 ^ mul_34_17_n_10931);
 assign mul_34_17_n_10421 = ~((mul_34_17_n_10904 | mul_34_17_n_10900) & (mul_34_17_n_10902 | mul_34_17_n_10901));
 assign mul_34_17_n_10420 = ~(mul_34_17_n_10361 & mul_34_17_n_10347);
 assign mul_34_17_n_10419 = ~(mul_34_17_n_10393 & mul_34_17_n_10352);
 assign mul_34_17_n_10418 = (mul_34_17_n_10861 ^ mul_34_17_n_10870);
 assign mul_34_17_n_10417 = (mul_34_17_n_10867 ^ mul_34_17_n_10860);
 assign mul_34_17_n_10416 = ~(mul_34_17_n_10348 | mul_34_17_n_10346);
 assign mul_34_17_n_10415 = ~mul_34_17_n_10375;
 assign mul_34_17_n_10414 = ~mul_34_17_n_10374;
 assign mul_34_17_n_10410 = ~mul_34_17_n_10409;
 assign mul_34_17_n_10408 = ~mul_34_17_n_10372;
 assign mul_34_17_n_10404 = ~mul_34_17_n_10405;
 assign mul_34_17_n_10400 = ~mul_34_17_n_10401;
 assign mul_34_17_n_10393 = ~mul_34_17_n_10394;
 assign mul_34_17_n_10391 = ~mul_34_17_n_10390;
 assign mul_34_17_n_10389 = ~mul_34_17_n_10388;
 assign mul_34_17_n_10383 = ~mul_34_17_n_10384;
 assign mul_34_17_n_10381 = ~mul_34_17_n_10380;
 assign mul_34_17_n_10377 = ~mul_34_17_n_10376;
 assign mul_34_17_n_10375 = ~(mul_34_17_n_11006 | mul_34_17_n_11000);
 assign mul_34_17_n_10374 = ~(mul_34_17_n_11046 | mul_34_17_n_11041);
 assign mul_34_17_n_10413 = ~(mul_34_17_n_10830 | mul_34_17_n_10884);
 assign mul_34_17_n_10412 = ~(mul_34_17_n_11006 & mul_34_17_n_11000);
 assign mul_34_17_n_10373 = ~(mul_34_17_n_10971 | mul_34_17_n_11251);
 assign mul_34_17_n_10411 = ~(mul_34_17_n_10877 | mul_34_17_n_10903);
 assign mul_34_17_n_10409 = ~(mul_34_17_n_10839 | mul_34_17_n_10881);
 assign mul_34_17_n_10372 = ~(mul_34_17_n_10951 | mul_34_17_n_10918);
 assign mul_34_17_n_10407 = ~(mul_34_17_n_10864 | mul_34_17_n_10841);
 assign mul_34_17_n_10406 = ~(mul_34_17_n_11016 | mul_34_17_n_10832);
 assign mul_34_17_n_10371 = ~(mul_34_17_n_10831 & mul_34_17_n_11024);
 assign mul_34_17_n_10405 = ~(mul_34_17_n_10924 & mul_34_17_n_10922);
 assign mul_34_17_n_10370 = ~(mul_34_17_n_10867 | mul_34_17_n_10860);
 assign mul_34_17_n_10403 = ~(mul_34_17_n_10967 | mul_34_17_n_10970);
 assign mul_34_17_n_10402 = ~(mul_34_17_n_10868 & mul_34_17_n_11030);
 assign mul_34_17_n_10401 = ~(mul_34_17_n_10983 & mul_34_17_n_10946);
 assign mul_34_17_n_10399 = ~(mul_34_17_n_11004 & mul_34_17_n_11050);
 assign mul_34_17_n_10398 = ~(mul_34_17_n_10944 | mul_34_17_n_10949);
 assign mul_34_17_n_10397 = ~(mul_34_17_n_10867 & mul_34_17_n_10860);
 assign mul_34_17_n_10396 = ~(mul_34_17_n_10838 | mul_34_17_n_10926);
 assign mul_34_17_n_10369 = ~(mul_34_17_n_10875 | mul_34_17_n_11019);
 assign mul_34_17_n_10395 = ~(mul_34_17_n_10887 & mul_34_17_n_10888);
 assign mul_34_17_n_10394 = ~(mul_34_17_n_10844 | mul_34_17_n_10966);
 assign mul_34_17_n_10392 = ~(mul_34_17_n_10880 | mul_34_17_n_10878);
 assign mul_34_17_n_10390 = ~(mul_34_17_n_10939 & mul_34_17_n_10931);
 assign mul_34_17_n_10368 = ~(mul_34_17_n_10827 | mul_34_17_n_10893);
 assign mul_34_17_n_10388 = ~(mul_34_17_n_10847 | mul_34_17_n_10886);
 assign mul_34_17_n_10387 = ~(mul_34_17_n_11003 & mul_34_17_n_10849);
 assign mul_34_17_n_10367 = ~(mul_34_17_n_10827 & mul_34_17_n_10893);
 assign mul_34_17_n_10386 = ~(mul_34_17_n_10902 | mul_34_17_n_10901);
 assign mul_34_17_n_10385 = ~(mul_34_17_n_11023 | mul_34_17_n_10879);
 assign mul_34_17_n_10384 = ~(mul_34_17_n_11046 | mul_34_17_n_10942);
 assign mul_34_17_n_10382 = ~(mul_34_17_n_10997 | mul_34_17_n_10828);
 assign mul_34_17_n_10380 = ~(mul_34_17_n_10944 & mul_34_17_n_10949);
 assign mul_34_17_n_10379 = ~(mul_34_17_n_10904 | mul_34_17_n_10900);
 assign mul_34_17_n_10378 = ~(mul_34_17_n_10876 | mul_34_17_n_11017);
 assign mul_34_17_n_10376 = ~(mul_34_17_n_10964 & mul_34_17_n_11011);
 assign mul_34_17_n_10366 = ~mul_34_17_n_10328;
 assign mul_34_17_n_10362 = ~mul_34_17_n_10363;
 assign mul_34_17_n_10356 = ~mul_34_17_n_10355;
 assign mul_34_17_n_10354 = ~mul_34_17_n_10353;
 assign mul_34_17_n_10350 = ~mul_34_17_n_10349;
 assign mul_34_17_n_10346 = ~mul_34_17_n_10347;
 assign mul_34_17_n_10345 = ~mul_34_17_n_10344;
 assign mul_34_17_n_10342 = ~mul_34_17_n_10343;
 assign mul_34_17_n_10340 = ~mul_34_17_n_10341;
 assign mul_34_17_n_10338 = ~mul_34_17_n_10339;
 assign mul_34_17_n_10337 = ~(mul_34_17_n_10836 | mul_34_17_n_10287);
 assign mul_34_17_n_10336 = ~(mul_34_17_n_10866 | mul_34_17_n_10930);
 assign mul_34_17_n_10335 = ~(mul_34_17_n_10295 & mul_34_17_n_11248);
 assign mul_34_17_n_10334 = ~(mul_34_17_n_11046 | mul_34_17_n_10299);
 assign mul_34_17_n_10333 = ~(mul_34_17_n_10294 & mul_34_17_n_10972);
 assign mul_34_17_n_10332 = ~(mul_34_17_n_11038 | mul_34_17_n_10292);
 assign mul_34_17_n_10331 = ~(mul_34_17_n_10999 | mul_34_17_n_11020);
 assign mul_34_17_n_10330 = ~(mul_34_17_n_10872 | mul_34_17_n_10312);
 assign mul_34_17_n_10329 = ~(mul_34_17_n_10942 | mul_34_17_n_10310);
 assign mul_34_17_n_10328 = ~(mul_34_17_n_10829 | mul_34_17_n_11047);
 assign mul_34_17_n_10327 = ~(mul_34_17_n_10967 | mul_34_17_n_10318);
 assign mul_34_17_n_10326 = ~(mul_34_17_n_10923 | mul_34_17_n_11031);
 assign mul_34_17_n_10325 = ~(mul_34_17_n_10881 | mul_34_17_n_10309);
 assign mul_34_17_n_10365 = ~(mul_34_17_n_10998 & mul_34_17_n_10899);
 assign mul_34_17_n_10324 = ~(mul_34_17_n_11022 | mul_34_17_n_10307);
 assign mul_34_17_n_10323 = ~(mul_34_17_n_10908 | mul_34_17_n_10286);
 assign mul_34_17_n_10322 = ~(mul_34_17_n_10947 & mul_34_17_n_10948);
 assign mul_34_17_n_10364 = ~(mul_34_17_n_10848 & mul_34_17_n_11025);
 assign mul_34_17_n_10321 = ~(mul_34_17_n_10940 | mul_34_17_n_10300);
 assign mul_34_17_n_10320 = ~(mul_34_17_n_10864 | mul_34_17_n_10296);
 assign mul_34_17_n_10363 = ~(mul_34_17_n_10955 | mul_34_17_n_10995);
 assign mul_34_17_n_10361 = ~(mul_34_17_n_11007 & mul_34_17_n_10842);
 assign mul_34_17_n_10360 = ~(mul_34_17_n_10850 | mul_34_17_n_11002);
 assign mul_34_17_n_10359 = ~(mul_34_17_n_10907 | mul_34_17_n_11018);
 assign mul_34_17_n_10358 = ~(mul_34_17_n_10941 | mul_34_17_n_10316);
 assign mul_34_17_n_10357 = ~(mul_34_17_n_10885 & mul_34_17_n_10856);
 assign mul_34_17_n_10355 = ~(mul_34_17_n_10876 & mul_34_17_n_11017);
 assign mul_34_17_n_10353 = ~(mul_34_17_n_10952 | mul_34_17_n_10911);
 assign mul_34_17_n_10352 = ~(mul_34_17_n_10844 & mul_34_17_n_10966);
 assign mul_34_17_n_10351 = ~(mul_34_17_n_10951 & mul_34_17_n_10918);
 assign mul_34_17_n_10349 = ~(mul_34_17_n_10896 & mul_34_17_n_10897);
 assign mul_34_17_n_10348 = ~(mul_34_17_n_10859 | mul_34_17_n_10858);
 assign mul_34_17_n_10347 = ~(mul_34_17_n_10859 & mul_34_17_n_10858);
 assign mul_34_17_n_10344 = ~(mul_34_17_n_10896 | mul_34_17_n_10897);
 assign mul_34_17_n_10343 = ~(mul_34_17_n_10829 & mul_34_17_n_11047);
 assign mul_34_17_n_10341 = ~(mul_34_17_n_10952 & mul_34_17_n_10911);
 assign mul_34_17_n_10339 = ~(mul_34_17_n_10887 | mul_34_17_n_10888);
 assign mul_34_17_n_10319 = ~mul_34_17_n_10933;
 assign mul_34_17_n_10318 = ~mul_34_17_n_10969;
 assign mul_34_17_n_10317 = ~mul_34_17_n_10866;
 assign mul_34_17_n_10316 = ~mul_34_17_n_10940;
 assign mul_34_17_n_10315 = ~mul_34_17_n_10826;
 assign mul_34_17_n_10314 = ~mul_34_17_n_10972;
 assign mul_34_17_n_10313 = ~mul_34_17_n_11247;
 assign mul_34_17_n_10312 = ~mul_34_17_n_11035;
 assign mul_34_17_n_10311 = ~mul_34_17_n_11252;
 assign mul_34_17_n_10310 = ~mul_34_17_n_11041;
 assign mul_34_17_n_10309 = ~mul_34_17_n_10883;
 assign mul_34_17_n_10308 = ~mul_34_17_n_10993;
 assign mul_34_17_n_10307 = ~mul_34_17_n_10882;
 assign mul_34_17_n_10306 = ~mul_34_17_n_10942;
 assign mul_34_17_n_10305 = ~mul_34_17_n_10872;
 assign mul_34_17_n_10304 = ~mul_34_17_n_11038;
 assign mul_34_17_n_10303 = ~mul_34_17_n_11024;
 assign mul_34_17_n_10302 = ~mul_34_17_n_10914;
 assign mul_34_17_n_10301 = ~mul_34_17_n_10845;
 assign mul_34_17_n_10300 = ~mul_34_17_n_10941;
 assign mul_34_17_n_10299 = ~mul_34_17_n_10912;
 assign mul_34_17_n_10298 = ~mul_34_17_n_10994;
 assign mul_34_17_n_10297 = ~mul_34_17_n_10953;
 assign mul_34_17_n_10296 = ~mul_34_17_n_11034;
 assign mul_34_17_n_10295 = ~mul_34_17_n_10864;
 assign mul_34_17_n_10294 = ~mul_34_17_n_10971;
 assign mul_34_17_n_10293 = ~mul_34_17_n_10831;
 assign mul_34_17_n_10292 = ~mul_34_17_n_10843;
 assign mul_34_17_n_10291 = ~mul_34_17_n_11022;
 assign mul_34_17_n_10290 = ~mul_34_17_n_10881;
 assign mul_34_17_n_10289 = ~mul_34_17_n_10890;
 assign mul_34_17_n_10288 = ~mul_34_17_n_10908;
 assign mul_34_17_n_10287 = ~mul_34_17_n_11042;
 assign mul_34_17_n_10286 = ~mul_34_17_n_10909;
 assign asc001_68_ = (mul_34_17_n_10790 ^ mul_34_17_n_10585);
 assign mul_34_17_n_10284 = ~mul_34_17_n_10285;
 assign mul_34_17_n_10285 = ~(mul_34_17_n_10774 & mul_34_17_n_10673);
 assign mul_34_17_n_10282 = ~mul_34_17_n_10283;
 assign mul_34_17_n_10283 = ~(mul_34_17_n_10437 & mul_34_17_n_10365);
 assign mul_34_17_n_10281 = ~(mul_34_17_n_10171 | mul_34_17_n_10270);
 assign mul_34_17_n_10280 = ~(mul_34_17_n_10245 & mul_34_17_n_10246);
 assign mul_34_17_n_10279 = ~(mul_34_17_n_10244 & mul_34_17_n_10247);
 assign mul_34_17_n_10278 = ((mul_34_17_n_10133 & mul_34_17_n_10185) | (mul_34_17_n_10229 & mul_34_17_n_10228));
 assign mul_34_17_n_10277 = ~(mul_34_17_n_10253 & mul_34_17_n_10254);
 assign mul_34_17_n_10276 = ~(mul_34_17_n_10251 & mul_34_17_n_10217);
 assign mul_34_17_n_10275 = ~(mul_34_17_n_10252 | mul_34_17_n_10216);
 assign mul_34_17_n_10274 = ~(mul_34_17_n_10004 & mul_34_17_n_10249);
 assign mul_34_17_n_10273 = ~(mul_34_17_n_10005 & mul_34_17_n_10250);
 assign mul_34_17_n_10272 = ~(mul_34_17_n_10219 | mul_34_17_n_338);
 assign mul_34_17_n_10271 = ~mul_34_17_n_10270;
 assign mul_34_17_n_10269 = ((mul_34_17_n_10082 & mul_34_17_n_10012) | ((mul_34_17_n_10082 & mul_34_17_n_10160)
    | (mul_34_17_n_10160 & mul_34_17_n_10012)));
 assign mul_34_17_n_10268 = ~(mul_34_17_n_10243 | mul_34_17_n_339);
 assign mul_34_17_n_10267 = ~(mul_34_17_n_10082 & mul_34_17_n_10248);
 assign mul_34_17_n_10266 = ~(mul_34_17_n_10253 | mul_34_17_n_10254);
 assign mul_34_17_n_10265 = ~(mul_34_17_n_10219 & mul_34_17_n_338);
 assign mul_34_17_n_10264 = ~(mul_34_17_n_10251 | mul_34_17_n_10217);
 assign mul_34_17_n_10263 = ~(mul_34_17_n_9959 ^ mul_34_17_n_10190);
 assign mul_34_17_n_10262 = ~(mul_34_17_n_9994 ^ mul_34_17_n_10189);
 assign mul_34_17_n_10261 = ~(mul_34_17_n_10193 ^ mul_34_17_n_10003);
 assign mul_34_17_n_10260 = ~(mul_34_17_n_10007 ^ mul_34_17_n_10192);
 assign mul_34_17_n_10259 = ~(mul_34_17_n_10194 ^ mul_34_17_n_10031);
 assign mul_34_17_n_10258 = ~(mul_34_17_n_10139 ^ mul_34_17_n_10187);
 assign mul_34_17_n_10270 = ~(mul_34_17_n_11286 ^ mul_34_17_n_10188);
 assign mul_34_17_n_10257 = ~(mul_34_17_n_10220 | mul_34_17_n_10215);
 assign mul_34_17_n_10256 = ~(mul_34_17_n_10220 & mul_34_17_n_10215);
 assign mul_34_17_n_10255 = ~(mul_34_17_n_9995 | mul_34_17_n_10214);
 assign mul_34_17_n_10250 = ~mul_34_17_n_10249;
 assign mul_34_17_n_10247 = ~mul_34_17_n_10246;
 assign mul_34_17_n_10245 = ~mul_34_17_n_10244;
 assign mul_34_17_n_10242 = ((mul_34_17_n_10108 & mul_34_17_n_10099) | ((mul_34_17_n_10108 & mul_34_17_n_10058)
    | (mul_34_17_n_10058 & mul_34_17_n_10099)));
 assign mul_34_17_n_10241 = ~(mul_34_17_n_10100 | mul_34_17_n_10218);
 assign mul_34_17_n_10240 = ~(mul_34_17_n_10100 & mul_34_17_n_10218);
 assign mul_34_17_n_10239 = ((mul_34_17_n_9990 & mul_34_17_n_9860) | (mul_34_17_n_10156 & mul_34_17_n_9955));
 assign mul_34_17_n_10238 = ((mul_34_17_n_9931 & mul_34_17_n_10027) | (mul_34_17_n_9913 & mul_34_17_n_10154));
 assign mul_34_17_n_10237 = ((mul_34_17_n_11276 & mul_34_17_n_10096) | ((mul_34_17_n_11276 & mul_34_17_n_10083)
    | (mul_34_17_n_10083 & mul_34_17_n_10096)));
 assign mul_34_17_n_10236 = ((mul_34_17_n_10086 & mul_34_17_n_10055) | ((mul_34_17_n_10086 & mul_34_17_n_9991)
    | (mul_34_17_n_9991 & mul_34_17_n_10055)));
 assign mul_34_17_n_10235 = ~(mul_34_17_n_10176 ^ mul_34_17_n_9888);
 assign mul_34_17_n_10234 = ~(mul_34_17_n_10158 ^ mul_34_17_n_332);
 assign mul_34_17_n_10233 = ~(mul_34_17_n_10157 ^ mul_34_17_n_9955);
 assign mul_34_17_n_10254 = ~(mul_34_17_n_10142 ^ mul_34_17_n_10006);
 assign mul_34_17_n_10253 = ((mul_34_17_n_11286 & mul_34_17_n_9961) | ((mul_34_17_n_11286 & mul_34_17_n_10088)
    | (mul_34_17_n_10088 & mul_34_17_n_9961)));
 assign mul_34_17_n_10252 = ((mul_34_17_n_9735 & mul_34_17_n_10020) | ((mul_34_17_n_9735 & mul_34_17_n_10102)
    | (mul_34_17_n_10102 & mul_34_17_n_10020)));
 assign mul_34_17_n_10251 = ~(mul_34_17_n_11278 ^ mul_34_17_n_10174);
 assign mul_34_17_n_10249 = ~(mul_34_17_n_10162 ^ mul_34_17_n_11284);
 assign mul_34_17_n_10248 = (mul_34_17_n_10160 ^ mul_34_17_n_10012);
 assign mul_34_17_n_10246 = ((mul_34_17_n_9999 & mul_34_17_n_10008) | ((mul_34_17_n_9999 & mul_34_17_n_10085)
    | (mul_34_17_n_10085 & mul_34_17_n_10008)));
 assign mul_34_17_n_10244 = ~((mul_34_17_n_9707 & (~mul_34_17_n_9908 & ~mul_34_17_n_10140)) | ((mul_34_17_n_9706
    & (mul_34_17_n_9908 & ~mul_34_17_n_10140)) | (mul_34_17_n_10087 & mul_34_17_n_10140)));
 assign mul_34_17_n_10243 = ((mul_34_17_n_10005 & mul_34_17_n_10163) | ((mul_34_17_n_10005 & mul_34_17_n_11284)
    | (mul_34_17_n_11284 & mul_34_17_n_10163)));
 assign mul_34_17_n_10232 = ~(mul_34_17_n_10108 ^ mul_34_17_n_10058);
 assign mul_34_17_n_10231 = ~(mul_34_17_n_10157 & mul_34_17_n_9954);
 assign mul_34_17_n_10230 = ~(mul_34_17_n_10161 | mul_34_17_n_10164);
 assign mul_34_17_n_10229 = ~(mul_34_17_n_10159 & mul_34_17_n_332);
 assign mul_34_17_n_10228 = ~(mul_34_17_n_10158 & mul_34_17_n_10081);
 assign mul_34_17_n_10227 = ~(mul_34_17_n_10134 & (mul_34_17_n_10135 & (mul_34_17_n_9974 & mul_34_17_n_9886)));
 assign mul_34_17_n_10226 = ~(mul_34_17_n_10094 & mul_34_17_n_10165);
 assign mul_34_17_n_10225 = ~(mul_34_17_n_9958 | mul_34_17_n_10166);
 assign mul_34_17_n_10224 = ~(mul_34_17_n_10172 | mul_34_17_n_10084);
 assign mul_34_17_n_10223 = ~(mul_34_17_n_9735 ^ mul_34_17_n_10102);
 assign mul_34_17_n_10222 = ~(mul_34_17_n_10042 & mul_34_17_n_10144);
 assign mul_34_17_n_10221 = ~(mul_34_17_n_9770 | (mul_34_17_n_10039 | (mul_34_17_n_9629 | mul_34_17_n_10123)));
 assign mul_34_17_n_10213 = ~(mul_34_17_n_9957 | mul_34_17_n_10167);
 assign mul_34_17_n_10212 = ((mul_34_17_n_9850 & mul_34_17_n_9943) | (mul_34_17_n_10107 & mul_34_17_n_9929));
 assign mul_34_17_n_10211 = ~(mul_34_17_n_10103 ^ mul_34_17_n_9932);
 assign mul_34_17_n_10210 = ~(mul_34_17_n_10168 | mul_34_17_n_9950);
 assign mul_34_17_n_10209 = ((mul_34_17_n_10093 & mul_34_17_n_9959) | (mul_34_17_n_9947 & mul_34_17_n_10051));
 assign mul_34_17_n_10208 = ((mul_34_17_n_317 & mul_34_17_n_11278) | ((mul_34_17_n_317 & mul_34_17_n_10029)
    | (mul_34_17_n_10029 & mul_34_17_n_11278)));
 assign mul_34_17_n_10207 = ((mul_34_17_n_10019 & mul_34_17_n_10033) | ((mul_34_17_n_10019 & mul_34_17_n_9737)
    | (mul_34_17_n_9737 & mul_34_17_n_10033)));
 assign mul_34_17_n_10206 = ~((mul_34_17_n_9931 | mul_34_17_n_10027) & (mul_34_17_n_10090 | mul_34_17_n_9913));
 assign mul_34_17_n_10205 = ~(mul_34_17_n_10061 ^ mul_34_17_n_9874);
 assign mul_34_17_n_10204 = ~(mul_34_17_n_10173 | mul_34_17_n_10085);
 assign mul_34_17_n_10203 = ~(mul_34_17_n_11282 ^ mul_34_17_n_10095);
 assign mul_34_17_n_10202 = ~(mul_34_17_n_9849 ^ mul_34_17_n_10066);
 assign mul_34_17_n_10201 = ((mul_34_17_n_10007 & mul_34_17_n_10060) | ((mul_34_17_n_10007 & mul_34_17_n_9977)
    | (mul_34_17_n_9977 & mul_34_17_n_10060)));
 assign mul_34_17_n_10200 = ((mul_34_17_n_10000 & mul_34_17_n_10098) | ((mul_34_17_n_10000 & mul_34_17_n_9779)
    | (mul_34_17_n_9779 & mul_34_17_n_10098)));
 assign mul_34_17_n_10199 = ~(mul_34_17_n_10065 ^ mul_34_17_n_9933);
 assign mul_34_17_n_10198 = ~(mul_34_17_n_10063 ^ mul_34_17_n_9871);
 assign mul_34_17_n_10197 = ~(mul_34_17_n_11306 ^ mul_34_17_n_10062);
 assign mul_34_17_n_10196 = ((mul_34_17_n_11274 & mul_34_17_n_332) | ((mul_34_17_n_11274 & mul_34_17_n_9996)
    | (mul_34_17_n_9996 & mul_34_17_n_332)));
 assign mul_34_17_n_10195 = ((mul_34_17_n_9584 & mul_34_17_n_10021) | ((mul_34_17_n_9584 & mul_34_17_n_9993)
    | (mul_34_17_n_9993 & mul_34_17_n_10021)));
 assign mul_34_17_n_10194 = ~(mul_34_17_n_10106 ^ mul_34_17_n_9928);
 assign mul_34_17_n_10193 = ~(mul_34_17_n_10089 ^ mul_34_17_n_10001);
 assign mul_34_17_n_10220 = ((mul_34_17_n_9976 & mul_34_17_n_9957) | ((mul_34_17_n_9976 & mul_34_17_n_9800)
    | (mul_34_17_n_9800 & mul_34_17_n_9957)));
 assign mul_34_17_n_10219 = ((mul_34_17_n_10002 & mul_34_17_n_10089) | ((mul_34_17_n_10002 & mul_34_17_n_10003)
    | (mul_34_17_n_10003 & mul_34_17_n_10089)));
 assign mul_34_17_n_10192 = ~(mul_34_17_n_9841 ^ (mul_34_17_n_9828 ^ (mul_34_17_n_9344 ^ mul_34_17_n_9927)));
 assign mul_34_17_n_10191 = (mul_34_17_n_11276 ^ mul_34_17_n_10096);
 assign mul_34_17_n_10190 = ~(mul_34_17_n_10059 ^ mul_34_17_n_10092);
 assign mul_34_17_n_10189 = ~(mul_34_17_n_9879 ^ (mul_34_17_n_9971 ^ (mul_34_17_n_9357 ^ mul_34_17_n_9625)));
 assign mul_34_17_n_10218 = ~((mul_34_17_n_9818 & (~mul_34_17_n_9906 & ~mul_34_17_n_10010)) | ((mul_34_17_n_9819
    & (mul_34_17_n_9906 & ~mul_34_17_n_10010)) | (mul_34_17_n_10071 & mul_34_17_n_10010)));
 assign mul_34_17_n_10188 = ~(mul_34_17_n_9961 ^ mul_34_17_n_10088);
 assign mul_34_17_n_10217 = ((mul_34_17_n_9997 & mul_34_17_n_10097) | ((mul_34_17_n_9997 & mul_34_17_n_11617)
    | (mul_34_17_n_11617 & mul_34_17_n_10097)));
 assign mul_34_17_n_10187 = ~(mul_34_17_n_9695 ^ mul_34_17_n_11272);
 assign mul_34_17_n_10216 = ~(mul_34_17_n_10009 ^ mul_34_17_n_10068);
 assign mul_34_17_n_10215 = ~(mul_34_17_n_9821 ^ (mul_34_17_n_9953 ^ (mul_34_17_n_9884 ^ mul_34_17_n_9725)));
 assign mul_34_17_n_10214 = ~(mul_34_17_n_11288 ^ mul_34_17_n_10067);
 assign mul_34_17_n_10186 = ~(mul_34_17_n_10111 & mul_34_17_n_10101);
 assign mul_34_17_n_10185 = ~(mul_34_17_n_10087 & mul_34_17_n_10114);
 assign mul_34_17_n_10184 = ~(mul_34_17_n_9931 ^ mul_34_17_n_10027);
 assign mul_34_17_n_10183 = ~((mul_34_17_n_9885 & mul_34_17_n_9797) | (mul_34_17_n_9847 & mul_34_17_n_10023));
 assign mul_34_17_n_10182 = ~(mul_34_17_n_10104 | mul_34_17_n_10109);
 assign mul_34_17_n_10181 = ~(mul_34_17_n_10111 | mul_34_17_n_10101);
 assign mul_34_17_n_10180 = ~(mul_34_17_n_10016 | mul_34_17_n_322);
 assign mul_34_17_n_10179 = ~(mul_34_17_n_10016 & mul_34_17_n_322);
 assign mul_34_17_n_10178 = ~((mul_34_17_n_10019 | mul_34_17_n_9737) & (mul_34_17_n_9833 | mul_34_17_n_9918));
 assign mul_34_17_n_10177 = ~(mul_34_17_n_10019 ^ mul_34_17_n_9737);
 assign mul_34_17_n_10176 = ~(mul_34_17_n_9847 ^ mul_34_17_n_10023);
 assign mul_34_17_n_10175 = ~(mul_34_17_n_10103 | mul_34_17_n_9932);
 assign mul_34_17_n_10174 = (mul_34_17_n_317 ^ mul_34_17_n_10029);
 assign mul_34_17_n_10173 = ~mul_34_17_n_10172;
 assign mul_34_17_n_10171 = ~mul_34_17_n_10170;
 assign mul_34_17_n_10169 = ~mul_34_17_n_10168;
 assign mul_34_17_n_10167 = ~mul_34_17_n_10166;
 assign mul_34_17_n_10163 = ~mul_34_17_n_10162;
 assign mul_34_17_n_10159 = ~mul_34_17_n_10158;
 assign mul_34_17_n_10156 = ~mul_34_17_n_10157;
 assign mul_34_17_n_10155 = ((mul_34_17_n_9909 & mul_34_17_n_9917) | ((mul_34_17_n_9909 & mul_34_17_n_9817)
    | (mul_34_17_n_9817 & mul_34_17_n_9917)));
 assign mul_34_17_n_10154 = ~(mul_34_17_n_10091 | mul_34_17_n_10112);
 assign mul_34_17_n_10153 = ((mul_34_17_n_9794 & mul_34_17_n_10035) | ((mul_34_17_n_9794 & mul_34_17_n_9926)
    | (mul_34_17_n_9926 & mul_34_17_n_10035)));
 assign mul_34_17_n_10152 = ~((mul_34_17_n_9764 & mul_34_17_n_9765) | (mul_34_17_n_10006 & mul_34_17_n_9998));
 assign mul_34_17_n_10151 = ((mul_34_17_n_10054 | mul_34_17_n_9968) & (mul_34_17_n_9479 | mul_34_17_n_9537));
 assign mul_34_17_n_10150 = ~(mul_34_17_n_10050 | mul_34_17_n_10095);
 assign mul_34_17_n_10149 = ((mul_34_17_n_9994 | mul_34_17_n_9799) & (mul_34_17_n_10048 | mul_34_17_n_10047));
 assign mul_34_17_n_10148 = ((mul_34_17_n_318 & mul_34_17_n_11304) | ((mul_34_17_n_318 & mul_34_17_n_9720)
    | (mul_34_17_n_9720 & mul_34_17_n_11304)));
 assign mul_34_17_n_10147 = ((mul_34_17_n_9887 & mul_34_17_n_9979) | ((mul_34_17_n_9887 & mul_34_17_n_9951)
    | (mul_34_17_n_9951 & mul_34_17_n_9979)));
 assign mul_34_17_n_10146 = ((mul_34_17_n_9712 & mul_34_17_n_10009) | ((mul_34_17_n_9712 & mul_34_17_n_9910)
    | (mul_34_17_n_9910 & mul_34_17_n_10009)));
 assign mul_34_17_n_10145 = (mul_34_17_n_9993 ^ mul_34_17_n_9584);
 assign mul_34_17_n_10144 = ((mul_34_17_n_9911 | mul_34_17_n_9709) & (mul_34_17_n_11288 | mul_34_17_n_9995));
 assign mul_34_17_n_10143 = ~((mul_34_17_n_9670 & mul_34_17_n_9964) | (mul_34_17_n_9969 & mul_34_17_n_10057));
 assign mul_34_17_n_10142 = ~(mul_34_17_n_9429 ^ (mul_34_17_n_9621 ^ (mul_34_17_n_9881 ^ mul_34_17_n_9727)));
 assign mul_34_17_n_10141 = ((mul_34_17_n_9866 & mul_34_17_n_9758) | (mul_34_17_n_333 & mul_34_17_n_10044));
 assign mul_34_17_n_10172 = (mul_34_17_n_9999 ^ mul_34_17_n_10008);
 assign mul_34_17_n_10140 = ~(mul_34_17_n_10055 ^ mul_34_17_n_9991);
 assign mul_34_17_n_10170 = ((mul_34_17_n_9953 & mul_34_17_n_9978) | ((mul_34_17_n_9953 & mul_34_17_n_9821)
    | (mul_34_17_n_9821 & mul_34_17_n_9978)));
 assign mul_34_17_n_10139 = ((mul_34_17_n_9787 & mul_34_17_n_10011) | ((mul_34_17_n_9787 & mul_34_17_n_9815)
    | (mul_34_17_n_9815 & mul_34_17_n_10011)));
 assign mul_34_17_n_10138 = (mul_34_17_n_9997 ^ mul_34_17_n_11617);
 assign mul_34_17_n_10168 = ~(mul_34_17_n_9732 ^ (mul_34_17_n_9882 ^ (mul_34_17_n_9286 ^ mul_34_17_n_9740)));
 assign mul_34_17_n_10137 = ~(mul_34_17_n_9774 ^ mul_34_17_n_10026);
 assign mul_34_17_n_10136 = ~(mul_34_17_n_10000 ^ mul_34_17_n_9779);
 assign mul_34_17_n_10166 = ~(mul_34_17_n_9846 ^ (mul_34_17_n_11296 ^ (mul_34_17_n_9213 ^ mul_34_17_n_9626)));
 assign mul_34_17_n_10165 = ~(mul_34_17_n_9982 ^ mul_34_17_n_9791);
 assign mul_34_17_n_10164 = ~(mul_34_17_n_10130 & mul_34_17_n_10052);
 assign mul_34_17_n_10162 = ~(mul_34_17_n_9785 ^ mul_34_17_n_9981);
 assign mul_34_17_n_10161 = ~(mul_34_17_n_9983 ^ mul_34_17_n_10011);
 assign mul_34_17_n_10160 = ~(mul_34_17_n_9880 ^ mul_34_17_n_9980);
 assign mul_34_17_n_10158 = (mul_34_17_n_11274 ^ mul_34_17_n_9996);
 assign mul_34_17_n_10157 = ((mul_34_17_n_9986 & mul_34_17_n_9902) | (mul_34_17_n_10046 & mul_34_17_n_9930));
 assign mul_34_17_n_10135 = ~(mul_34_17_n_9773 & mul_34_17_n_10025);
 assign mul_34_17_n_10134 = ~(mul_34_17_n_9774 & mul_34_17_n_10026);
 assign mul_34_17_n_10133 = ~(mul_34_17_n_9985 & mul_34_17_n_9992);
 assign mul_34_17_n_10132 = ~(mul_34_17_n_10015 | mul_34_17_n_10024);
 assign mul_34_17_n_10131 = ~(mul_34_17_n_9794 ^ mul_34_17_n_9926);
 assign mul_34_17_n_10130 = ((mul_34_17_n_9768 & mul_34_17_n_9868) | (mul_34_17_n_9889 & mul_34_17_n_9783));
 assign mul_34_17_n_10129 = ~(mul_34_17_n_10006 | mul_34_17_n_9998);
 assign mul_34_17_n_10128 = ~(mul_34_17_n_10036 | mul_34_17_n_10010);
 assign mul_34_17_n_10127 = ~(mul_34_17_n_10015 & mul_34_17_n_10024);
 assign mul_34_17_n_10126 = ~(mul_34_17_n_9870 | mul_34_17_n_10013);
 assign mul_34_17_n_10125 = ~(mul_34_17_n_9869 | mul_34_17_n_10014);
 assign mul_34_17_n_10124 = ~(mul_34_17_n_9872 | mul_34_17_n_10017);
 assign mul_34_17_n_10123 = ~(mul_34_17_n_10054 | mul_34_17_n_9966);
 assign mul_34_17_n_10122 = ~(mul_34_17_n_11288 & mul_34_17_n_9995);
 assign mul_34_17_n_10121 = ~(mul_34_17_n_9873 | mul_34_17_n_10018);
 assign mul_34_17_n_10120 = ~((mul_34_17_n_9761 & mul_34_17_n_9763) | (mul_34_17_n_9945 & mul_34_17_n_9861));
 assign mul_34_17_n_10119 = ~(mul_34_17_n_9877 & (mul_34_17_n_9561 & (mul_34_17_n_9795 & mul_34_17_n_9967)));
 assign mul_34_17_n_10118 = ~(mul_34_17_n_9729 ^ mul_34_17_n_303);
 assign mul_34_17_n_10117 = (mul_34_17_n_9833 ^ mul_34_17_n_9918);
 assign mul_34_17_n_10116 = ~(mul_34_17_n_10054 & mul_34_17_n_10056);
 assign mul_34_17_n_10115 = ~(mul_34_17_n_9811 & mul_34_17_n_10028);
 assign mul_34_17_n_10114 = ~(mul_34_17_n_10055 & mul_34_17_n_9991);
 assign mul_34_17_n_10113 = ~(mul_34_17_n_9847 | mul_34_17_n_10023);
 assign mul_34_17_n_10112 = ~(mul_34_17_n_9931 | mul_34_17_n_10027);
 assign mul_34_17_n_10110 = ~mul_34_17_n_10109;
 assign mul_34_17_n_10107 = ~mul_34_17_n_10106;
 assign mul_34_17_n_10105 = ~mul_34_17_n_10104;
 assign mul_34_17_n_10093 = ~mul_34_17_n_10092;
 assign mul_34_17_n_10091 = ~mul_34_17_n_10090;
 assign mul_34_17_n_10087 = ~mul_34_17_n_10086;
 assign mul_34_17_n_10084 = ~mul_34_17_n_10085;
 assign mul_34_17_n_10081 = ~mul_34_17_n_332;
 assign mul_34_17_n_10080 = ~((mul_34_17_n_9631 & mul_34_17_n_9760) | (mul_34_17_n_9776 & mul_34_17_n_300));
 assign mul_34_17_n_10079 = ((mul_34_17_n_9739 & mul_34_17_n_9972) | ((mul_34_17_n_9739 & mul_34_17_n_9682)
    | (mul_34_17_n_9682 & mul_34_17_n_9972)));
 assign mul_34_17_n_10078 = ((mul_34_17_n_11292 & mul_34_17_n_9962) | ((mul_34_17_n_11292 & mul_34_17_n_9843)
    | (mul_34_17_n_9843 & mul_34_17_n_9962)));
 assign mul_34_17_n_10077 = ((mul_34_17_n_9715 & mul_34_17_n_9916) | ((mul_34_17_n_9715 & mul_34_17_n_9874)
    | (mul_34_17_n_9874 & mul_34_17_n_9916)));
 assign mul_34_17_n_10076 = ((mul_34_17_n_9778 & mul_34_17_n_9924) | ((mul_34_17_n_9778 & mul_34_17_n_11306)
    | (mul_34_17_n_11306 & mul_34_17_n_9924)));
 assign mul_34_17_n_10075 = ~(mul_34_17_n_9891 ^ mul_34_17_n_9690);
 assign mul_34_17_n_10074 = ~(mul_34_17_n_9920 ^ mul_34_17_n_9895);
 assign mul_34_17_n_10073 = ((mul_34_17_n_9274 & mul_34_17_n_9921) | ((mul_34_17_n_9274 & mul_34_17_n_9713)
    | (mul_34_17_n_9713 & mul_34_17_n_9921)));
 assign mul_34_17_n_10072 = ((mul_34_17_n_9689 & mul_34_17_n_9791) | ((mul_34_17_n_9689 & mul_34_17_n_9798)
    | (mul_34_17_n_9798 & mul_34_17_n_9791)));
 assign mul_34_17_n_10071 = ~(mul_34_17_n_9906 ^ mul_34_17_n_9818);
 assign mul_34_17_n_10111 = ~(mul_34_17_n_9921 ^ mul_34_17_n_9898);
 assign mul_34_17_n_10109 = ((mul_34_17_n_9822 & mul_34_17_n_11298) | ((mul_34_17_n_9822 & mul_34_17_n_9869)
    | (mul_34_17_n_9869 & mul_34_17_n_11298)));
 assign mul_34_17_n_10108 = ~(mul_34_17_n_9936 ^ mul_34_17_n_9832);
 assign mul_34_17_n_10106 = ~(mul_34_17_n_9973 ^ mul_34_17_n_9825);
 assign mul_34_17_n_10069 = ((mul_34_17_n_9593 & mul_34_17_n_9920) | ((mul_34_17_n_9593 & mul_34_17_n_9719)
    | (mul_34_17_n_9719 & mul_34_17_n_9920)));
 assign mul_34_17_n_10104 = ~(mul_34_17_n_9896 ^ mul_34_17_n_9837);
 assign mul_34_17_n_10103 = ~(mul_34_17_n_9549 ^ mul_34_17_n_9900);
 assign mul_34_17_n_10068 = (mul_34_17_n_9910 ^ mul_34_17_n_9712);
 assign mul_34_17_n_10102 = ~(mul_34_17_n_11310 ^ mul_34_17_n_9894);
 assign mul_34_17_n_10067 = (mul_34_17_n_9911 ^ mul_34_17_n_9709);
 assign mul_34_17_n_10101 = ((mul_34_17_n_9816 & mul_34_17_n_9366) | ((mul_34_17_n_9816 & mul_34_17_n_9773)
    | (mul_34_17_n_9773 & mul_34_17_n_9366)));
 assign mul_34_17_n_10066 = ~(mul_34_17_n_9775 ^ mul_34_17_n_300);
 assign mul_34_17_n_10065 = ~(mul_34_17_n_9772 ^ (mul_34_17_n_9782 ^ (mul_34_17_n_9099 ^ mul_34_17_n_9553)));
 assign mul_34_17_n_10064 = (mul_34_17_n_9917 ^ mul_34_17_n_9817);
 assign mul_34_17_n_10063 = ~(mul_34_17_n_306 ^ (mul_34_17_n_9726 ^ (mul_34_17_n_9300 ^ mul_34_17_n_9504)));
 assign mul_34_17_n_10062 = ~(mul_34_17_n_9777 ^ mul_34_17_n_9923);
 assign mul_34_17_n_10061 = ~(mul_34_17_n_9714 ^ mul_34_17_n_9915);
 assign mul_34_17_n_10100 = ((mul_34_17_n_9871 & mul_34_17_n_9890) | ((mul_34_17_n_9871 & mul_34_17_n_9687)
    | (mul_34_17_n_9687 & mul_34_17_n_9890)));
 assign mul_34_17_n_10099 = ((mul_34_17_n_9583 & mul_34_17_n_9930) | ((mul_34_17_n_9583 & mul_34_17_n_9820)
    | (mul_34_17_n_9820 & mul_34_17_n_9930)));
 assign mul_34_17_n_10060 = ~(mul_34_17_n_9344 ^ mul_34_17_n_9927);
 assign mul_34_17_n_10098 = ((mul_34_17_n_9807 & mul_34_17_n_9840) | (mul_34_17_n_9903 & mul_34_17_n_9755));
 assign mul_34_17_n_10097 = ((mul_34_17_n_9611 & mul_34_17_n_9922) | ((mul_34_17_n_9611 & mul_34_17_n_9616)
    | (mul_34_17_n_9616 & mul_34_17_n_9922)));
 assign mul_34_17_n_10096 = ~(mul_34_17_n_351 ^ mul_34_17_n_9937);
 assign mul_34_17_n_10095 = ~(mul_34_17_n_9901 ^ mul_34_17_n_9468);
 assign mul_34_17_n_10094 = ((mul_34_17_n_9873 & mul_34_17_n_9835) | ((mul_34_17_n_9873 & mul_34_17_n_9585)
    | (mul_34_17_n_9585 & mul_34_17_n_9835)));
 assign mul_34_17_n_10092 = ~(mul_34_17_n_318 ^ mul_34_17_n_9907);
 assign mul_34_17_n_10090 = ~(mul_34_17_n_9892 ^ mul_34_17_n_9654);
 assign mul_34_17_n_10059 = ((mul_34_17_n_9880 & mul_34_17_n_9975) | (mul_34_17_n_291 & mul_34_17_n_9590));
 assign mul_34_17_n_10089 = ~(mul_34_17_n_9922 ^ mul_34_17_n_9854);
 assign mul_34_17_n_10088 = ~(mul_34_17_n_11300 ^ mul_34_17_n_9893);
 assign mul_34_17_n_10086 = ~(mul_34_17_n_9908 ^ mul_34_17_n_9706);
 assign mul_34_17_n_10085 = ~(mul_34_17_n_9899 ^ mul_34_17_n_9789);
 assign mul_34_17_n_10083 = ((mul_34_17_n_9663 & mul_34_17_n_9960) | ((mul_34_17_n_9663 & mul_34_17_n_9780)
    | (mul_34_17_n_9780 & mul_34_17_n_9960)));
 assign mul_34_17_n_10082 = ((mul_34_17_n_9591 & mul_34_17_n_9827) | ((mul_34_17_n_9591 & mul_34_17_n_9811)
    | (mul_34_17_n_9811 & mul_34_17_n_9827)));
 assign mul_34_17_n_10057 = ~mul_34_17_n_10056;
 assign mul_34_17_n_10053 = ~(mul_34_17_n_9679 & mul_34_17_n_9925);
 assign mul_34_17_n_10052 = ~(mul_34_17_n_9948 & mul_34_17_n_9784);
 assign mul_34_17_n_10051 = ~(mul_34_17_n_9880 & mul_34_17_n_9975);
 assign mul_34_17_n_10050 = ~(mul_34_17_n_9914 | mul_34_17_n_11282);
 assign mul_34_17_n_10049 = ~(mul_34_17_n_318 & mul_34_17_n_9907);
 assign mul_34_17_n_10048 = ~(mul_34_17_n_9879 | mul_34_17_n_9970);
 assign mul_34_17_n_10047 = ~(mul_34_17_n_9878 | mul_34_17_n_9971);
 assign mul_34_17_n_10046 = ~(mul_34_17_n_9583 ^ mul_34_17_n_9820);
 assign mul_34_17_n_10045 = ~(mul_34_17_n_9776 | mul_34_17_n_300);
 assign mul_34_17_n_10044 = ~(mul_34_17_n_9973 & mul_34_17_n_9825);
 assign mul_34_17_n_10043 = ~(mul_34_17_n_9845 ^ mul_34_17_n_11302);
 assign mul_34_17_n_10042 = ~(mul_34_17_n_9911 & mul_34_17_n_9709);
 assign mul_34_17_n_10041 = ~(mul_34_17_n_11292 ^ mul_34_17_n_9843);
 assign mul_34_17_n_10040 = ~(mul_34_17_n_9679 | mul_34_17_n_9925);
 assign mul_34_17_n_10039 = ~(mul_34_17_n_9747 | mul_34_17_n_9965);
 assign mul_34_17_n_10038 = ((mul_34_17_n_11292 & mul_34_17_n_9843) | (mul_34_17_n_9844 & mul_34_17_n_9612));
 assign mul_34_17_n_10037 = ~(mul_34_17_n_9818 | mul_34_17_n_9906);
 assign mul_34_17_n_10036 = ~(mul_34_17_n_9819 | mul_34_17_n_9905);
 assign mul_34_17_n_10058 = ((mul_34_17_n_350 & mul_34_17_n_9559) | (mul_34_17_n_9863 & mul_34_17_n_9406));
 assign mul_34_17_n_10035 = ~(mul_34_17_n_9729 & mul_34_17_n_303);
 assign mul_34_17_n_10034 = ~(mul_34_17_n_9974 & mul_34_17_n_9886);
 assign mul_34_17_n_10033 = ~(mul_34_17_n_9834 | mul_34_17_n_9919);
 assign mul_34_17_n_10032 = ~(mul_34_17_n_9833 | mul_34_17_n_9918);
 assign mul_34_17_n_10056 = ~(mul_34_17_n_9877 & (mul_34_17_n_9561 & (mul_34_17_n_9684 & mul_34_17_n_301)));
 assign mul_34_17_n_10031 = ((mul_34_17_n_9678 & mul_34_17_n_351) | ((mul_34_17_n_9678 & mul_34_17_n_294)
    | (mul_34_17_n_294 & mul_34_17_n_351)));
 assign mul_34_17_n_10055 = ((mul_34_17_n_352 & mul_34_17_n_9789) | ((mul_34_17_n_352 & mul_34_17_n_9660)
    | (mul_34_17_n_9660 & mul_34_17_n_9789)));
 assign mul_34_17_n_10030 = ~(mul_34_17_n_9794 & mul_34_17_n_9926);
 assign mul_34_17_n_10054 = ~(mul_34_17_n_9752 | mul_34_17_n_9940);
 assign mul_34_17_n_10025 = ~mul_34_17_n_10026;
 assign mul_34_17_n_10022 = ~mul_34_17_n_10021;
 assign mul_34_17_n_10018 = ~mul_34_17_n_10017;
 assign mul_34_17_n_10014 = ~mul_34_17_n_10013;
 assign mul_34_17_n_10004 = ~mul_34_17_n_10005;
 assign mul_34_17_n_10002 = ~mul_34_17_n_10001;
 assign mul_34_17_n_9992 = ~mul_34_17_n_9991;
 assign mul_34_17_n_9990 = ~(mul_34_17_n_9859 & mul_34_17_n_9920);
 assign mul_34_17_n_9989 = ((mul_34_17_n_236 & mul_34_17_n_9877) | ((mul_34_17_n_236 & mul_34_17_n_8791)
    | (mul_34_17_n_8791 & mul_34_17_n_9877)));
 assign mul_34_17_n_9988 = ~(mul_34_17_n_9802 ^ mul_34_17_n_9601);
 assign mul_34_17_n_9987 = ((mul_34_17_n_9743 & mul_34_17_n_9825) | ((mul_34_17_n_9743 & mul_34_17_n_9609)
    | (mul_34_17_n_9609 & mul_34_17_n_9825)));
 assign mul_34_17_n_9986 = (mul_34_17_n_9583 ^ mul_34_17_n_9820);
 assign mul_34_17_n_9985 = ((mul_34_17_n_9385 & mul_34_17_n_9867) | (mul_34_17_n_9851 & mul_34_17_n_11290));
 assign mul_34_17_n_9984 = ((mul_34_17_n_9686 & mul_34_17_n_9549) | ((mul_34_17_n_9686 & mul_34_17_n_9445)
    | (mul_34_17_n_9445 & mul_34_17_n_9549)));
 assign mul_34_17_n_10029 = ((mul_34_17_n_287 & mul_34_17_n_9836) | ((mul_34_17_n_287 & mul_34_17_n_9542)
    | (mul_34_17_n_9542 & mul_34_17_n_9836)));
 assign mul_34_17_n_9983 = (mul_34_17_n_9787 ^ mul_34_17_n_9815);
 assign mul_34_17_n_10028 = (mul_34_17_n_9591 ^ mul_34_17_n_9827);
 assign mul_34_17_n_10027 = ~(mul_34_17_n_11280 ^ mul_34_17_n_9697);
 assign mul_34_17_n_10026 = (mul_34_17_n_9816 ^ mul_34_17_n_9366);
 assign mul_34_17_n_10024 = ~(mul_34_17_n_9790 ^ mul_34_17_n_9805);
 assign mul_34_17_n_9982 = ~(mul_34_17_n_8987 ^ (mul_34_17_n_9498 ^ (mul_34_17_n_9547 ^ mul_34_17_n_9614)));
 assign mul_34_17_n_10023 = ~(mul_34_17_n_9801 ^ mul_34_17_n_9831);
 assign mul_34_17_n_9981 = ~(mul_34_17_n_9587 ^ mul_34_17_n_9829);
 assign mul_34_17_n_10021 = ((mul_34_17_n_9788 & mul_34_17_n_11312) | ((mul_34_17_n_9788 & mul_34_17_n_9475)
    | (mul_34_17_n_9475 & mul_34_17_n_11312)));
 assign mul_34_17_n_10020 = ((mul_34_17_n_9781 & mul_34_17_n_9490) | ((mul_34_17_n_9781 & mul_34_17_n_9468)
    | (mul_34_17_n_9468 & mul_34_17_n_9490)));
 assign mul_34_17_n_10019 = ~(mul_34_17_n_9853 ^ mul_34_17_n_9509);
 assign mul_34_17_n_9980 = ~(mul_34_17_n_9839 ^ mul_34_17_n_9590);
 assign mul_34_17_n_10017 = (mul_34_17_n_9585 ^ mul_34_17_n_9835);
 assign mul_34_17_n_10016 = ((mul_34_17_n_9722 & mul_34_17_n_9838) | ((mul_34_17_n_9722 & mul_34_17_n_9659)
    | (mul_34_17_n_9659 & mul_34_17_n_9838)));
 assign mul_34_17_n_10015 = ((mul_34_17_n_9532 & mul_34_17_n_11280) | ((mul_34_17_n_9532 & mul_34_17_n_9278)
    | (mul_34_17_n_9278 & mul_34_17_n_11280)));
 assign mul_34_17_n_10013 = (mul_34_17_n_11298 ^ mul_34_17_n_9822);
 assign mul_34_17_n_9979 = (mul_34_17_n_9732 ^ mul_34_17_n_9882);
 assign mul_34_17_n_10012 = ~((mul_34_17_n_299 & mul_34_17_n_9862) | (mul_34_17_n_9604 & mul_34_17_n_9809));
 assign mul_34_17_n_10011 = ((mul_34_17_n_9771 & mul_34_17_n_9489) | ((mul_34_17_n_9771 & mul_34_17_n_9426)
    | (mul_34_17_n_9426 & mul_34_17_n_9489)));
 assign mul_34_17_n_10010 = ~(mul_34_17_n_9602 ^ mul_34_17_n_9852);
 assign mul_34_17_n_9978 = (mul_34_17_n_9884 ^ mul_34_17_n_9725);
 assign mul_34_17_n_10009 = ((mul_34_17_n_9711 & mul_34_17_n_11310) | ((mul_34_17_n_9711 & mul_34_17_n_9473)
    | (mul_34_17_n_9473 & mul_34_17_n_11310)));
 assign mul_34_17_n_10008 = ((mul_34_17_n_9361 & mul_34_17_n_354) | (mul_34_17_n_9253 & mul_34_17_n_9864));
 assign mul_34_17_n_10007 = ((mul_34_17_n_9596 & mul_34_17_n_9840) | ((mul_34_17_n_9596 & mul_34_17_n_9595)
    | (mul_34_17_n_9595 & mul_34_17_n_9840)));
 assign mul_34_17_n_10006 = ((mul_34_17_n_9538 & mul_34_17_n_9672) | ((mul_34_17_n_9538 & mul_34_17_n_9710)
    | (mul_34_17_n_9710 & mul_34_17_n_9672)));
 assign mul_34_17_n_10005 = ((mul_34_17_n_9656 & mul_34_17_n_9708) | ((mul_34_17_n_9656 & mul_34_17_n_9721)
    | (mul_34_17_n_9721 & mul_34_17_n_9708)));
 assign mul_34_17_n_10003 = ((mul_34_17_n_9594 & mul_34_17_n_9828) | ((mul_34_17_n_9594 & mul_34_17_n_9599)
    | (mul_34_17_n_9599 & mul_34_17_n_9828)));
 assign mul_34_17_n_10001 = ~((mul_34_17_n_9702 & mul_34_17_n_9492) | (mul_34_17_n_9399 & mul_34_17_n_9858));
 assign mul_34_17_n_9977 = (mul_34_17_n_9841 ^ mul_34_17_n_9828);
 assign mul_34_17_n_10000 = ((mul_34_17_n_9786 & mul_34_17_n_9829) | ((mul_34_17_n_9786 & mul_34_17_n_9588)
    | (mul_34_17_n_9588 & mul_34_17_n_9829)));
 assign mul_34_17_n_9999 = ((mul_34_17_n_9655 & mul_34_17_n_9831) | ((mul_34_17_n_9655 & mul_34_17_n_9598)
    | (mul_34_17_n_9598 & mul_34_17_n_9831)));
 assign mul_34_17_n_9976 = (mul_34_17_n_9846 ^ mul_34_17_n_11296);
 assign mul_34_17_n_9998 = (mul_34_17_n_9881 ^ mul_34_17_n_9727);
 assign mul_34_17_n_9997 = ~(mul_34_17_n_9804 ^ mul_34_17_n_9836);
 assign mul_34_17_n_9996 = ((mul_34_17_n_9472 & mul_34_17_n_9724) | ((mul_34_17_n_9472 & mul_34_17_n_9706)
    | (mul_34_17_n_9706 & mul_34_17_n_9724)));
 assign mul_34_17_n_9995 = ((mul_34_17_n_9741 & mul_34_17_n_9879) | ((mul_34_17_n_9741 & mul_34_17_n_9619)
    | (mul_34_17_n_9619 & mul_34_17_n_9879)));
 assign mul_34_17_n_9994 = ((mul_34_17_n_11294 & mul_34_17_n_304) | (mul_34_17_n_9883 & mul_34_17_n_9832));
 assign mul_34_17_n_9993 = ~(mul_34_17_n_9803 ^ mul_34_17_n_9669);
 assign mul_34_17_n_9991 = ~(mul_34_17_n_11314 ^ mul_34_17_n_9806);
 assign mul_34_17_n_9970 = ~mul_34_17_n_9971;
 assign mul_34_17_n_9969 = ~mul_34_17_n_9968;
 assign mul_34_17_n_9967 = ~mul_34_17_n_9966;
 assign mul_34_17_n_9965 = ~mul_34_17_n_9964;
 assign mul_34_17_n_9963 = ~mul_34_17_n_9962;
 assign mul_34_17_n_9958 = ~mul_34_17_n_9957;
 assign mul_34_17_n_9955 = ~mul_34_17_n_9954;
 assign mul_34_17_n_9950 = ~mul_34_17_n_9951;
 assign mul_34_17_n_9949 = ~(mul_34_17_n_9830 | mul_34_17_n_9855);
 assign mul_34_17_n_9948 = ~(mul_34_17_n_9772 ^ mul_34_17_n_9782);
 assign mul_34_17_n_9947 = ~(mul_34_17_n_291 & mul_34_17_n_9590);
 assign mul_34_17_n_9975 = ~(mul_34_17_n_9839 & mul_34_17_n_9589);
 assign mul_34_17_n_9945 = ~(mul_34_17_n_9883 & mul_34_17_n_9832);
 assign mul_34_17_n_9943 = ~(mul_34_17_n_351 & mul_34_17_n_319);
 assign mul_34_17_n_9974 = ((mul_34_17_n_9391 & mul_34_17_n_9640) | (mul_34_17_n_9418 & mul_34_17_n_9734));
 assign mul_34_17_n_9942 = ~(mul_34_17_n_9793 | mul_34_17_n_9842);
 assign mul_34_17_n_9941 = ~(mul_34_17_n_9739 ^ mul_34_17_n_9682);
 assign mul_34_17_n_9940 = ((mul_34_17_n_9677 & mul_34_17_n_9795) | (mul_34_17_n_9376 & mul_34_17_n_9304));
 assign mul_34_17_n_9939 = ~(mul_34_17_n_9824 & mul_34_17_n_9823);
 assign mul_34_17_n_9938 = ~(mul_34_17_n_9824 | mul_34_17_n_9823);
 assign mul_34_17_n_9973 = ~(mul_34_17_n_9743 ^ mul_34_17_n_9609);
 assign mul_34_17_n_9972 = ~(mul_34_17_n_9793 & mul_34_17_n_9842);
 assign mul_34_17_n_9937 = ~(mul_34_17_n_9678 ^ mul_34_17_n_294);
 assign mul_34_17_n_9971 = (mul_34_17_n_9741 ^ mul_34_17_n_9619);
 assign mul_34_17_n_9936 = ~(mul_34_17_n_9606 ^ mul_34_17_n_9742);
 assign mul_34_17_n_9935 = ~(mul_34_17_n_9556 ^ mul_34_17_n_9792);
 assign mul_34_17_n_9968 = ~(mul_34_17_n_9670 & mul_34_17_n_9876);
 assign mul_34_17_n_9966 = ~(mul_34_17_n_305 & (mul_34_17_n_9670 & (mul_34_17_n_313 & mul_34_17_n_9543)));
 assign mul_34_17_n_9964 = ((mul_34_17_n_9369 & mul_34_17_n_9506) | ((mul_34_17_n_9369 & mul_34_17_n_9627)
    | (mul_34_17_n_9627 & mul_34_17_n_9506)));
 assign mul_34_17_n_9962 = ~(mul_34_17_n_9845 & mul_34_17_n_11302);
 assign mul_34_17_n_9934 = ~(mul_34_17_n_9844 & mul_34_17_n_9612);
 assign mul_34_17_n_9961 = ((mul_34_17_n_9618 & mul_34_17_n_9725) | ((mul_34_17_n_9618 & mul_34_17_n_9554)
    | (mul_34_17_n_9554 & mul_34_17_n_9725)));
 assign mul_34_17_n_9960 = ((mul_34_17_n_9177 & mul_34_17_n_11314) | ((mul_34_17_n_9177 & mul_34_17_n_9597)
    | (mul_34_17_n_9597 & mul_34_17_n_11314)));
 assign mul_34_17_n_9933 = ((mul_34_17_n_9658 & mul_34_17_n_9669) | ((mul_34_17_n_9658 & mul_34_17_n_9422)
    | (mul_34_17_n_9422 & mul_34_17_n_9669)));
 assign mul_34_17_n_9959 = ((mul_34_17_n_9530 & mul_34_17_n_9604) | ((mul_34_17_n_9530 & mul_34_17_n_9664)
    | (mul_34_17_n_9664 & mul_34_17_n_9604)));
 assign mul_34_17_n_9957 = ((mul_34_17_n_9375 & mul_34_17_n_9602) | ((mul_34_17_n_9375 & mul_34_17_n_9615)
    | (mul_34_17_n_9615 & mul_34_17_n_9602)));
 assign mul_34_17_n_9954 = ((mul_34_17_n_9662 & mul_34_17_n_9601) | ((mul_34_17_n_9662 & mul_34_17_n_9350)
    | (mul_34_17_n_9350 & mul_34_17_n_9601)));
 assign mul_34_17_n_9953 = ((mul_34_17_n_9533 & mul_34_17_n_9653) | ((mul_34_17_n_9533 & mul_34_17_n_9582)
    | (mul_34_17_n_9582 & mul_34_17_n_9653)));
 assign mul_34_17_n_9951 = ((mul_34_17_n_9558 & mul_34_17_n_9727) | ((mul_34_17_n_9558 & mul_34_17_n_9610)
    | (mul_34_17_n_9610 & mul_34_17_n_9727)));
 assign mul_34_17_n_9929 = ~mul_34_17_n_9928;
 assign mul_34_17_n_9924 = ~mul_34_17_n_9923;
 assign mul_34_17_n_9918 = ~mul_34_17_n_9919;
 assign mul_34_17_n_9916 = ~mul_34_17_n_9915;
 assign mul_34_17_n_9906 = ~mul_34_17_n_9905;
 assign mul_34_17_n_9903 = ~((mul_34_17_n_9581 & mul_34_17_n_9478) | (mul_34_17_n_309 & mul_34_17_n_9749));
 assign mul_34_17_n_9902 = ~(mul_34_17_n_9688 ^ mul_34_17_n_9463);
 assign mul_34_17_n_9901 = (mul_34_17_n_9781 ^ mul_34_17_n_9490);
 assign mul_34_17_n_9932 = ((mul_34_17_n_9661 & mul_34_17_n_9790) | ((mul_34_17_n_9661 & mul_34_17_n_9341)
    | (mul_34_17_n_9341 & mul_34_17_n_9790)));
 assign mul_34_17_n_9900 = ~(mul_34_17_n_9227 ^ (mul_34_17_n_9502 ^ (mul_34_17_n_9217 ^ mul_34_17_n_8859)));
 assign mul_34_17_n_9931 = ((mul_34_17_n_9654 & mul_34_17_n_9723) | ((mul_34_17_n_9654 & mul_34_17_n_9469)
    | (mul_34_17_n_9469 & mul_34_17_n_9723)));
 assign mul_34_17_n_9899 = (mul_34_17_n_352 ^ mul_34_17_n_9660);
 assign mul_34_17_n_9930 = ~(mul_34_17_n_9331 ^ (mul_34_17_n_9539 ^ (mul_34_17_n_9307 ^ mul_34_17_n_9092)));
 assign mul_34_17_n_9898 = (mul_34_17_n_9274 ^ mul_34_17_n_9713);
 assign mul_34_17_n_9897 = (mul_34_17_n_9663 ^ mul_34_17_n_9780);
 assign mul_34_17_n_9896 = (mul_34_17_n_9722 ^ mul_34_17_n_9659);
 assign mul_34_17_n_9895 = ~(mul_34_17_n_9118 ^ (mul_34_17_n_9373 ^ (mul_34_17_n_8927 ^ mul_34_17_n_9557)));
 assign mul_34_17_n_9928 = ((mul_34_17_n_353 & mul_34_17_n_9544) | (mul_34_17_n_9443 & mul_34_17_n_9796));
 assign mul_34_17_n_9894 = (mul_34_17_n_9711 ^ mul_34_17_n_9473);
 assign mul_34_17_n_9927 = ~(mul_34_17_n_9728 ^ mul_34_17_n_9343);
 assign mul_34_17_n_9926 = ~(mul_34_17_n_9179 ^ mul_34_17_n_9699);
 assign mul_34_17_n_9925 = ~(mul_34_17_n_9696 ^ mul_34_17_n_9419);
 assign mul_34_17_n_9893 = ~(mul_34_17_n_9710 ^ mul_34_17_n_9538);
 assign mul_34_17_n_9892 = ~(mul_34_17_n_9469 ^ mul_34_17_n_9723);
 assign mul_34_17_n_9891 = (mul_34_17_n_9734 ^ mul_34_17_n_9418);
 assign mul_34_17_n_9923 = ~(mul_34_17_n_9665 ^ mul_34_17_n_9746);
 assign mul_34_17_n_9922 = ((mul_34_17_n_9344 & mul_34_17_n_9728) | ((mul_34_17_n_9344 & mul_34_17_n_9343)
    | (mul_34_17_n_9343 & mul_34_17_n_9728)));
 assign mul_34_17_n_9921 = ~((mul_34_17_n_9117 & (~mul_34_17_n_9535 & ~mul_34_17_n_9430)) | ((mul_34_17_n_9116
    & (mul_34_17_n_9535 & ~mul_34_17_n_9430)) | (mul_34_17_n_9766 & mul_34_17_n_9430)));
 assign mul_34_17_n_9920 = ((mul_34_17_n_281 & mul_34_17_n_9733) | ((mul_34_17_n_281 & mul_34_17_n_9531)
    | (mul_34_17_n_9531 & mul_34_17_n_9733)));
 assign mul_34_17_n_9890 = (mul_34_17_n_306 ^ mul_34_17_n_9726);
 assign mul_34_17_n_9919 = ~(mul_34_17_n_9330 ^ mul_34_17_n_9693);
 assign mul_34_17_n_9917 = ~(mul_34_17_n_9694 ^ mul_34_17_n_9730);
 assign mul_34_17_n_9915 = ~(mul_34_17_n_9674 ^ mul_34_17_n_9748);
 assign mul_34_17_n_9914 = ((mul_34_17_n_9337 & mul_34_17_n_9730) | ((mul_34_17_n_9337 & mul_34_17_n_9476)
    | (mul_34_17_n_9476 & mul_34_17_n_9730)));
 assign mul_34_17_n_9889 = ~(mul_34_17_n_9771 ^ mul_34_17_n_9782);
 assign mul_34_17_n_9888 = ~(mul_34_17_n_9885 & mul_34_17_n_9797);
 assign mul_34_17_n_9913 = ((mul_34_17_n_9199 & mul_34_17_n_9570) | (mul_34_17_n_311 & mul_34_17_n_9392));
 assign mul_34_17_n_9887 = ~(mul_34_17_n_9286 ^ mul_34_17_n_9740);
 assign mul_34_17_n_9911 = ~(mul_34_17_n_9656 ^ mul_34_17_n_9721);
 assign mul_34_17_n_9910 = ~(mul_34_17_n_9700 ^ mul_34_17_n_9788);
 assign mul_34_17_n_9909 = ((mul_34_17_n_9481 & mul_34_17_n_9731) | ((mul_34_17_n_9481 & mul_34_17_n_9482)
    | (mul_34_17_n_9482 & mul_34_17_n_9731)));
 assign mul_34_17_n_9908 = (mul_34_17_n_9472 ^ mul_34_17_n_9724);
 assign mul_34_17_n_9907 = ~(mul_34_17_n_11304 ^ mul_34_17_n_9720);
 assign mul_34_17_n_9905 = ~((mul_34_17_n_9633 | mul_34_17_n_9726) & (mul_34_17_n_9365 | mul_34_17_n_9461));
 assign mul_34_17_n_9878 = ~mul_34_17_n_9879;
 assign mul_34_17_n_9876 = ~mul_34_17_n_9875;
 assign mul_34_17_n_9872 = ~mul_34_17_n_9873;
 assign mul_34_17_n_9870 = ~mul_34_17_n_9869;
 assign mul_34_17_n_9868 = ~(mul_34_17_n_9767 & mul_34_17_n_9669);
 assign mul_34_17_n_9867 = ~(mul_34_17_n_352 | mul_34_17_n_9514);
 assign mul_34_17_n_9886 = ~(mul_34_17_n_9417 & mul_34_17_n_308);
 assign mul_34_17_n_9885 = ((mul_34_17_n_9555 & mul_34_17_n_9666) | (mul_34_17_n_9522 & mul_34_17_n_9641));
 assign mul_34_17_n_9866 = ~(mul_34_17_n_9443 & mul_34_17_n_9796);
 assign mul_34_17_n_9865 = ~(mul_34_17_n_9605 & mul_34_17_n_9744);
 assign mul_34_17_n_9864 = ~(mul_34_17_n_9254 | mul_34_17_n_354);
 assign mul_34_17_n_9863 = ~(mul_34_17_n_350 | mul_34_17_n_9405);
 assign mul_34_17_n_9862 = ~(mul_34_17_n_9530 ^ mul_34_17_n_9664);
 assign mul_34_17_n_9861 = ~(mul_34_17_n_11294 & mul_34_17_n_304);
 assign mul_34_17_n_9860 = ~(mul_34_17_n_9593 & mul_34_17_n_9719);
 assign mul_34_17_n_9859 = ~(mul_34_17_n_9592 & mul_34_17_n_9718);
 assign mul_34_17_n_9858 = ~(mul_34_17_n_9703 | mul_34_17_n_9398);
 assign mul_34_17_n_9857 = ~(mul_34_17_n_9369 ^ mul_34_17_n_9627);
 assign mul_34_17_n_9856 = ~((mul_34_17_n_9511 & mul_34_17_n_9650) | (mul_34_17_n_9235 & mul_34_17_n_9409));
 assign mul_34_17_n_9855 = ~(mul_34_17_n_9556 | mul_34_17_n_9792);
 assign mul_34_17_n_9854 = ~(mul_34_17_n_9611 ^ mul_34_17_n_9616);
 assign mul_34_17_n_9853 = ~(mul_34_17_n_9199 ^ mul_34_17_n_9617);
 assign mul_34_17_n_9884 = ~(mul_34_17_n_9618 ^ mul_34_17_n_9554);
 assign mul_34_17_n_9852 = (mul_34_17_n_9375 ^ mul_34_17_n_9615);
 assign mul_34_17_n_9851 = ~(mul_34_17_n_352 & mul_34_17_n_9660);
 assign mul_34_17_n_9850 = ~(mul_34_17_n_9678 & mul_34_17_n_294);
 assign mul_34_17_n_9883 = ~(mul_34_17_n_9606 & mul_34_17_n_9742);
 assign mul_34_17_n_9882 = ~(mul_34_17_n_9555 ^ mul_34_17_n_9667);
 assign mul_34_17_n_9881 = ~(mul_34_17_n_9558 ^ mul_34_17_n_9610);
 assign mul_34_17_n_9880 = ((mul_34_17_n_279 & mul_34_17_n_9668) | ((mul_34_17_n_279 & mul_34_17_n_9440)
    | (mul_34_17_n_9440 & mul_34_17_n_9668)));
 assign mul_34_17_n_9879 = ((mul_34_17_n_283 & mul_34_17_n_9559) | ((mul_34_17_n_283 & mul_34_17_n_9480)
    | (mul_34_17_n_9480 & mul_34_17_n_9559)));
 assign mul_34_17_n_9877 = ~(mul_34_17_n_9757 & mul_34_17_n_9756);
 assign mul_34_17_n_9849 = ((mul_34_17_n_9535 & mul_34_17_n_9431) | ((mul_34_17_n_9535 & mul_34_17_n_9116)
    | (mul_34_17_n_9116 & mul_34_17_n_9431)));
 assign mul_34_17_n_9875 = ~((mul_34_17_n_9362 | mul_34_17_n_9438) & (mul_34_17_n_9369 | mul_34_17_n_9627));
 assign mul_34_17_n_9848 = ~(mul_34_17_n_9738 | mul_34_17_n_9681);
 assign mul_34_17_n_9874 = ((mul_34_17_n_9303 & mul_34_17_n_9665) | ((mul_34_17_n_9303 & mul_34_17_n_9497)
    | (mul_34_17_n_9497 & mul_34_17_n_9665)));
 assign mul_34_17_n_9873 = ((mul_34_17_n_9182 & mul_34_17_n_9600) | ((mul_34_17_n_9182 & mul_34_17_n_9342)
    | (mul_34_17_n_9342 & mul_34_17_n_9600)));
 assign mul_34_17_n_9871 = ((mul_34_17_n_9500 & mul_34_17_n_9674) | ((mul_34_17_n_9500 & mul_34_17_n_9439)
    | (mul_34_17_n_9439 & mul_34_17_n_9674)));
 assign mul_34_17_n_9869 = ((mul_34_17_n_9222 & mul_34_17_n_9359) | ((mul_34_17_n_9222 & mul_34_17_n_9503)
    | (mul_34_17_n_9503 & mul_34_17_n_9359)));
 assign mul_34_17_n_9844 = ~mul_34_17_n_9845;
 assign mul_34_17_n_9838 = ~mul_34_17_n_9837;
 assign mul_34_17_n_9833 = ~mul_34_17_n_9834;
 assign mul_34_17_n_9818 = ~mul_34_17_n_9819;
 assign mul_34_17_n_9809 = (mul_34_17_n_9664 ^ mul_34_17_n_9530);
 assign mul_34_17_n_9808 = ~(mul_34_17_n_9668 ^ mul_34_17_n_9637);
 assign mul_34_17_n_9807 = (mul_34_17_n_9596 ^ mul_34_17_n_9595);
 assign mul_34_17_n_9847 = ~(mul_34_17_n_9483 ^ mul_34_17_n_9568);
 assign mul_34_17_n_9846 = (mul_34_17_n_9533 ^ mul_34_17_n_9582);
 assign mul_34_17_n_9845 = ~(mul_34_17_n_9562 ^ mul_34_17_n_9271);
 assign mul_34_17_n_9806 = (mul_34_17_n_9177 ^ mul_34_17_n_9597);
 assign mul_34_17_n_9843 = ~(mul_34_17_n_9563 ^ mul_34_17_n_9283);
 assign mul_34_17_n_9842 = ~(mul_34_17_n_9567 ^ mul_34_17_n_9272);
 assign mul_34_17_n_9805 = ~(mul_34_17_n_9341 ^ mul_34_17_n_9661);
 assign mul_34_17_n_9804 = (mul_34_17_n_287 ^ mul_34_17_n_9542);
 assign mul_34_17_n_9803 = (mul_34_17_n_9658 ^ mul_34_17_n_9422);
 assign mul_34_17_n_9802 = (mul_34_17_n_9350 ^ mul_34_17_n_9662);
 assign mul_34_17_n_9841 = (mul_34_17_n_9594 ^ mul_34_17_n_9599);
 assign mul_34_17_n_9840 = ~(mul_34_17_n_9372 ^ (mul_34_17_n_8618 ^ (mul_34_17_n_9167 ^ mul_34_17_n_9174)));
 assign mul_34_17_n_9801 = (mul_34_17_n_9655 ^ mul_34_17_n_9598);
 assign mul_34_17_n_9839 = ~(mul_34_17_n_9423 ^ (mul_34_17_n_9296 ^ (mul_34_17_n_8952 ^ mul_34_17_n_8409)));
 assign mul_34_17_n_9837 = ~(mul_34_17_n_9546 ^ mul_34_17_n_9639);
 assign mul_34_17_n_9836 = ((mul_34_17_n_9492 & mul_34_17_n_9467) | ((mul_34_17_n_9492 & mul_34_17_n_9162)
    | (mul_34_17_n_9162 & mul_34_17_n_9467)));
 assign mul_34_17_n_9835 = ~(mul_34_17_n_9550 ^ mul_34_17_n_9634);
 assign mul_34_17_n_9834 = ((mul_34_17_n_9179 & mul_34_17_n_9491) | ((mul_34_17_n_9179 & mul_34_17_n_9540)
    | (mul_34_17_n_9540 & mul_34_17_n_9491)));
 assign mul_34_17_n_9832 = ((mul_34_17_n_9331 & mul_34_17_n_9463) | ((mul_34_17_n_9331 & mul_34_17_n_9539)
    | (mul_34_17_n_9539 & mul_34_17_n_9463)));
 assign mul_34_17_n_9831 = ((mul_34_17_n_9529 & mul_34_17_n_9286) | ((mul_34_17_n_9529 & mul_34_17_n_9336)
    | (mul_34_17_n_9336 & mul_34_17_n_9286)));
 assign mul_34_17_n_9830 = ~((mul_34_17_n_9182 & (~mul_34_17_n_9342 & ~mul_34_17_n_9600)) | ((mul_34_17_n_9181
    & (mul_34_17_n_9342 & ~mul_34_17_n_9600)) | (mul_34_17_n_9578 & mul_34_17_n_9600)));
 assign mul_34_17_n_9829 = ~((mul_34_17_n_357 & mul_34_17_n_9209) | (mul_34_17_n_9647 & mul_34_17_n_9078));
 assign mul_34_17_n_9828 = ((mul_34_17_n_9167 & mul_34_17_n_9581) | ((mul_34_17_n_9167 & mul_34_17_n_9175)
    | (mul_34_17_n_9175 & mul_34_17_n_9581)));
 assign mul_34_17_n_9827 = ((mul_34_17_n_9207 & mul_34_17_n_356) | (mul_34_17_n_9651 & mul_34_17_n_9084));
 assign mul_34_17_n_9825 = ((mul_34_17_n_9334 & mul_34_17_n_9485) | ((mul_34_17_n_9334 & mul_34_17_n_9470)
    | (mul_34_17_n_9470 & mul_34_17_n_9485)));
 assign mul_34_17_n_9800 = ~(mul_34_17_n_9213 ^ mul_34_17_n_9626);
 assign mul_34_17_n_9824 = ((mul_34_17_n_9419 & mul_34_17_n_8998) | (mul_34_17_n_9572 & mul_34_17_n_9393));
 assign mul_34_17_n_9823 = ~(mul_34_17_n_9566 ^ mul_34_17_n_9338);
 assign mul_34_17_n_9822 = ~(mul_34_17_n_9545 ^ mul_34_17_n_9569);
 assign mul_34_17_n_9821 = ~(mul_34_17_n_9295 ^ mul_34_17_n_9565);
 assign mul_34_17_n_9820 = ((mul_34_17_n_9268 & mul_34_17_n_9460) | (mul_34_17_n_9579 & mul_34_17_n_9082));
 assign mul_34_17_n_9819 = ~(mul_34_17_n_9191 ^ mul_34_17_n_9564);
 assign mul_34_17_n_9799 = (mul_34_17_n_9357 ^ mul_34_17_n_9625);
 assign mul_34_17_n_9798 = ~(mul_34_17_n_9547 ^ mul_34_17_n_9614);
 assign mul_34_17_n_9817 = ~(mul_34_17_n_9204 ^ mul_34_17_n_9632);
 assign mul_34_17_n_9816 = ~(mul_34_17_n_9638 ^ mul_34_17_n_9287);
 assign mul_34_17_n_9815 = ~(mul_34_17_n_9635 ^ mul_34_17_n_9551);
 assign mul_34_17_n_9811 = ((mul_34_17_n_9326 & mul_34_17_n_9411) | ((mul_34_17_n_9326 & mul_34_17_n_9544)
    | (mul_34_17_n_9544 & mul_34_17_n_9411)));
 assign mul_34_17_n_9786 = ~mul_34_17_n_9785;
 assign mul_34_17_n_9784 = ~mul_34_17_n_9783;
 assign mul_34_17_n_9778 = ~mul_34_17_n_9777;
 assign mul_34_17_n_9776 = ~mul_34_17_n_9775;
 assign mul_34_17_n_9773 = ~mul_34_17_n_9774;
 assign mul_34_17_n_9771 = ~mul_34_17_n_9772;
 assign mul_34_17_n_9770 = ~(mul_34_17_n_391 | mul_34_17_n_9636);
 assign mul_34_17_n_9768 = ~(mul_34_17_n_9658 & mul_34_17_n_9422);
 assign mul_34_17_n_9767 = ~(mul_34_17_n_9657 & mul_34_17_n_9421);
 assign mul_34_17_n_9766 = ~(mul_34_17_n_9535 ^ mul_34_17_n_9117);
 assign mul_34_17_n_9797 = ~(mul_34_17_n_11308 & mul_34_17_n_9667);
 assign mul_34_17_n_9765 = ~(mul_34_17_n_9429 & mul_34_17_n_9620);
 assign mul_34_17_n_9764 = ~(mul_34_17_n_9428 & mul_34_17_n_9621);
 assign mul_34_17_n_9763 = ~(mul_34_17_n_9357 & mul_34_17_n_9624);
 assign mul_34_17_n_9762 = ((mul_34_17_n_8855 & mul_34_17_n_9526) | ((mul_34_17_n_8855 & mul_34_17_n_8495)
    | (mul_34_17_n_8495 & mul_34_17_n_9526)));
 assign mul_34_17_n_9761 = ~(mul_34_17_n_11322 & mul_34_17_n_9625);
 assign mul_34_17_n_9760 = ~(mul_34_17_n_9431 & mul_34_17_n_9630);
 assign mul_34_17_n_9796 = ~(mul_34_17_n_353 | mul_34_17_n_9390);
 assign mul_34_17_n_9758 = ~(mul_34_17_n_353 & mul_34_17_n_9544);
 assign mul_34_17_n_9757 = ~(mul_34_17_n_9133 & mul_34_17_n_9675);
 assign mul_34_17_n_9756 = ~((mul_34_17_n_11334 & mul_34_17_n_8804) | (mul_34_17_n_9517 & mul_34_17_n_9526));
 assign mul_34_17_n_9755 = ~(mul_34_17_n_9580 & mul_34_17_n_9477);
 assign mul_34_17_n_9754 = ~(mul_34_17_n_9622 | mul_34_17_n_9608);
 assign mul_34_17_n_9753 = ~(mul_34_17_n_9441 & mul_34_17_n_9643);
 assign mul_34_17_n_9752 = ~(mul_34_17_n_9494 | mul_34_17_n_9646);
 assign mul_34_17_n_9751 = ~(mul_34_17_n_9374 ^ mul_34_17_n_9499);
 assign mul_34_17_n_9750 = ~(mul_34_17_n_9644 & mul_34_17_n_9676);
 assign mul_34_17_n_9795 = ((mul_34_17_n_9376 | mul_34_17_n_9304) & (mul_34_17_n_9495 | mul_34_17_n_9211));
 assign mul_34_17_n_9749 = ~(mul_34_17_n_9596 & mul_34_17_n_9595);
 assign mul_34_17_n_9748 = ~(mul_34_17_n_9500 ^ mul_34_17_n_9439);
 assign mul_34_17_n_9747 = ~(mul_34_17_n_305 & mul_34_17_n_9670);
 assign mul_34_17_n_9746 = (mul_34_17_n_9303 ^ mul_34_17_n_9497);
 assign mul_34_17_n_9794 = ((mul_34_17_n_9425 & mul_34_17_n_9548) | ((mul_34_17_n_9425 & mul_34_17_n_8990)
    | (mul_34_17_n_8990 & mul_34_17_n_9548)));
 assign mul_34_17_n_9793 = ((mul_34_17_n_9340 & mul_34_17_n_9301) | ((mul_34_17_n_9340 & mul_34_17_n_9283)
    | (mul_34_17_n_9283 & mul_34_17_n_9301)));
 assign mul_34_17_n_9792 = ((mul_34_17_n_9225 & mul_34_17_n_9546) | ((mul_34_17_n_9225 & mul_34_17_n_9370)
    | (mul_34_17_n_9370 & mul_34_17_n_9546)));
 assign mul_34_17_n_9745 = ~(mul_34_17_n_9222 ^ mul_34_17_n_9503);
 assign mul_34_17_n_9791 = ((mul_34_17_n_9220 & mul_34_17_n_9550) | ((mul_34_17_n_9220 & mul_34_17_n_9368)
    | (mul_34_17_n_9368 & mul_34_17_n_9550)));
 assign mul_34_17_n_9790 = ((mul_34_17_n_9094 & mul_34_17_n_355) | ((mul_34_17_n_9094 & mul_34_17_n_9100)
    | (mul_34_17_n_9100 & mul_34_17_n_355)));
 assign mul_34_17_n_9789 = ((mul_34_17_n_9333 & mul_34_17_n_9483) | ((mul_34_17_n_9333 & mul_34_17_n_9196)
    | (mul_34_17_n_9196 & mul_34_17_n_9483)));
 assign mul_34_17_n_9744 = ~(mul_34_17_n_9530 & mul_34_17_n_9664);
 assign mul_34_17_n_9788 = ((mul_34_17_n_9223 & mul_34_17_n_9447) | ((mul_34_17_n_9223 & mul_34_17_n_9037)
    | (mul_34_17_n_9037 & mul_34_17_n_9447)));
 assign mul_34_17_n_9787 = ((mul_34_17_n_9435 & mul_34_17_n_9402) | (mul_34_17_n_9519 & mul_34_17_n_9257));
 assign mul_34_17_n_9785 = ((mul_34_17_n_9356 & mul_34_17_n_9493) | ((mul_34_17_n_9356 & mul_34_17_n_11316)
    | (mul_34_17_n_11316 & mul_34_17_n_9493)));
 assign mul_34_17_n_9783 = ~(mul_34_17_n_9099 ^ mul_34_17_n_9553);
 assign mul_34_17_n_9782 = ~(mul_34_17_n_9426 ^ mul_34_17_n_9489);
 assign mul_34_17_n_9781 = ((mul_34_17_n_9228 & mul_34_17_n_9204) | ((mul_34_17_n_9228 & mul_34_17_n_277)
    | (mul_34_17_n_277 & mul_34_17_n_9204)));
 assign mul_34_17_n_9780 = ~(mul_34_17_n_9134 ^ mul_34_17_n_9512);
 assign mul_34_17_n_9779 = ((mul_34_17_n_9354 & mul_34_17_n_276) | ((mul_34_17_n_9354 & mul_34_17_n_9352)
    | (mul_34_17_n_9352 & mul_34_17_n_276)));
 assign mul_34_17_n_9777 = ((mul_34_17_n_9415 & mul_34_17_n_9547) | ((mul_34_17_n_9415 & mul_34_17_n_9180)
    | (mul_34_17_n_9180 & mul_34_17_n_9547)));
 assign mul_34_17_n_9775 = ((mul_34_17_n_358 & mul_34_17_n_9046) | (mul_34_17_n_9520 & mul_34_17_n_8911));
 assign mul_34_17_n_9774 = ((mul_34_17_n_282 & mul_34_17_n_9527) | ((mul_34_17_n_282 & mul_34_17_n_9120)
    | (mul_34_17_n_9120 & mul_34_17_n_9527)));
 assign mul_34_17_n_9772 = ((mul_34_17_n_9433 & mul_34_17_n_9130) | ((mul_34_17_n_9433 & mul_34_17_n_8929)
    | (mul_34_17_n_8929 & mul_34_17_n_9130)));
 assign mul_34_17_n_9739 = ~mul_34_17_n_9738;
 assign mul_34_17_n_9719 = ~mul_34_17_n_9718;
 assign mul_34_17_n_9715 = ~mul_34_17_n_9714;
 assign mul_34_17_n_9708 = ~mul_34_17_n_9709;
 assign mul_34_17_n_9707 = ~mul_34_17_n_9706;
 assign mul_34_17_n_9704 = (mul_34_17_n_9479 ^ mul_34_17_n_9537);
 assign mul_34_17_n_9703 = (mul_34_17_n_9467 ^ mul_34_17_n_9162);
 assign mul_34_17_n_9702 = (mul_34_17_n_9162 ^ mul_34_17_n_9467);
 assign mul_34_17_n_9700 = ~(mul_34_17_n_11312 ^ mul_34_17_n_9475);
 assign mul_34_17_n_9743 = ~(mul_34_17_n_9451 ^ mul_34_17_n_9093);
 assign mul_34_17_n_9699 = ~(mul_34_17_n_9491 ^ mul_34_17_n_9540);
 assign mul_34_17_n_9698 = ~(mul_34_17_n_9548 ^ mul_34_17_n_8990);
 assign mul_34_17_n_9742 = ~(mul_34_17_n_9262 ^ mul_34_17_n_9474);
 assign mul_34_17_n_9697 = ~(mul_34_17_n_9532 ^ mul_34_17_n_9278);
 assign mul_34_17_n_9696 = ~(mul_34_17_n_9455 ^ mul_34_17_n_8831);
 assign mul_34_17_n_9741 = ~(mul_34_17_n_9202 ^ mul_34_17_n_9507);
 assign mul_34_17_n_9740 = ~(mul_34_17_n_9529 ^ mul_34_17_n_9336);
 assign mul_34_17_n_9738 = ~(mul_34_17_n_9434 ^ mul_34_17_n_9450);
 assign mul_34_17_n_9695 = ((mul_34_17_n_9424 & mul_34_17_n_9552) | ((mul_34_17_n_9424 & mul_34_17_n_9420)
    | (mul_34_17_n_9420 & mul_34_17_n_9552)));
 assign mul_34_17_n_9694 = (mul_34_17_n_9337 ^ mul_34_17_n_9476);
 assign mul_34_17_n_9693 = ~(mul_34_17_n_9042 ^ (mul_34_17_n_8375 ^ (mul_34_17_n_9229 ^ mul_34_17_n_9297)));
 assign mul_34_17_n_9737 = ((mul_34_17_n_9330 & mul_34_17_n_9446) | ((mul_34_17_n_9330 & mul_34_17_n_9309)
    | (mul_34_17_n_9309 & mul_34_17_n_9446)));
 assign mul_34_17_n_9692 = (mul_34_17_n_9482 ^ mul_34_17_n_9481);
 assign mul_34_17_n_9691 = (mul_34_17_n_281 ^ mul_34_17_n_9531);
 assign mul_34_17_n_9735 = ((mul_34_17_n_9172 & mul_34_17_n_9166) | ((mul_34_17_n_9172 & mul_34_17_n_9325)
    | (mul_34_17_n_9325 & mul_34_17_n_9166)));
 assign mul_34_17_n_9690 = ((mul_34_17_n_9560 & mul_34_17_n_8953) | (mul_34_17_n_271 & mul_34_17_n_9105));
 assign mul_34_17_n_9734 = ~(mul_34_17_n_9536 ^ mul_34_17_n_9527);
 assign mul_34_17_n_9733 = ((mul_34_17_n_9423 & mul_34_17_n_9296) | ((mul_34_17_n_9423 & mul_34_17_n_9159)
    | (mul_34_17_n_9159 & mul_34_17_n_9296)));
 assign mul_34_17_n_9732 = ((mul_34_17_n_9349 & mul_34_17_n_9429) | ((mul_34_17_n_9349 & mul_34_17_n_9282)
    | (mul_34_17_n_9282 & mul_34_17_n_9429)));
 assign mul_34_17_n_9731 = ((mul_34_17_n_9189 & mul_34_17_n_9329) | ((mul_34_17_n_9189 & mul_34_17_n_9328)
    | (mul_34_17_n_9328 & mul_34_17_n_9329)));
 assign mul_34_17_n_9730 = ((mul_34_17_n_9160 & mul_34_17_n_9466) | ((mul_34_17_n_9160 & mul_34_17_n_9332)
    | (mul_34_17_n_9332 & mul_34_17_n_9466)));
 assign mul_34_17_n_9729 = ((mul_34_17_n_9339 & mul_34_17_n_290) | ((mul_34_17_n_9339 & mul_34_17_n_9187)
    | (mul_34_17_n_9187 & mul_34_17_n_290)));
 assign mul_34_17_n_9728 = ~((mul_34_17_n_8602 & (~mul_34_17_n_9164 & ~mul_34_17_n_8637)) | ((mul_34_17_n_8601
    & (mul_34_17_n_9164 & ~mul_34_17_n_8637)) | (mul_34_17_n_9458 & mul_34_17_n_8637)));
 assign mul_34_17_n_9727 = ((mul_34_17_n_9158 & mul_34_17_n_11320) | ((mul_34_17_n_9158 & mul_34_17_n_286)
    | (mul_34_17_n_286 & mul_34_17_n_11320)));
 assign mul_34_17_n_9726 = ((mul_34_17_n_9346 & mul_34_17_n_9239) | ((mul_34_17_n_9346 & mul_34_17_n_266)
    | (mul_34_17_n_266 & mul_34_17_n_9239)));
 assign mul_34_17_n_9725 = ((mul_34_17_n_9193 & mul_34_17_n_9213) | ((mul_34_17_n_9193 & mul_34_17_n_280)
    | (mul_34_17_n_280 & mul_34_17_n_9213)));
 assign mul_34_17_n_9724 = ((mul_34_17_n_9327 & mul_34_17_n_9462) | ((mul_34_17_n_9327 & mul_34_17_n_9361)
    | (mul_34_17_n_9361 & mul_34_17_n_9462)));
 assign mul_34_17_n_9723 = ~(mul_34_17_n_9448 ^ mul_34_17_n_9121);
 assign mul_34_17_n_9722 = ((mul_34_17_n_9188 & mul_34_17_n_9545) | ((mul_34_17_n_9188 & mul_34_17_n_9353)
    | (mul_34_17_n_9353 & mul_34_17_n_9545)));
 assign mul_34_17_n_9721 = ~(mul_34_17_n_9000 ^ mul_34_17_n_9452);
 assign mul_34_17_n_9689 = (mul_34_17_n_8987 ^ mul_34_17_n_9498);
 assign mul_34_17_n_9720 = ~(mul_34_17_n_11326 ^ mul_34_17_n_9513);
 assign mul_34_17_n_9718 = (mul_34_17_n_8927 ^ mul_34_17_n_9557);
 assign mul_34_17_n_9688 = (mul_34_17_n_9331 ^ mul_34_17_n_9539);
 assign mul_34_17_n_9717 = ((mul_34_17_n_9436 & mul_34_17_n_8986) | ((mul_34_17_n_9436 & mul_34_17_n_8913)
    | (mul_34_17_n_8913 & mul_34_17_n_8986)));
 assign mul_34_17_n_9716 = ~((mul_34_17_n_8543 & (~mul_34_17_n_0 & ~mul_34_17_n_9505)) | ((mul_34_17_n_8544
    & (mul_34_17_n_0 & ~mul_34_17_n_9505)) | (mul_34_17_n_9524 & mul_34_17_n_9505)));
 assign mul_34_17_n_9687 = ~(mul_34_17_n_9300 ^ mul_34_17_n_9504);
 assign mul_34_17_n_9714 = ~((mul_34_17_n_266 & (~mul_34_17_n_9284 & ~mul_34_17_n_9347)) | ((mul_34_17_n_8828
    & (mul_34_17_n_9284 & ~mul_34_17_n_9347)) | (mul_34_17_n_9457 & mul_34_17_n_9347)));
 assign mul_34_17_n_9686 = (mul_34_17_n_9227 ^ mul_34_17_n_9502);
 assign mul_34_17_n_9713 = ((mul_34_17_n_9115 & mul_34_17_n_9287) | ((mul_34_17_n_9115 & mul_34_17_n_9416)
    | (mul_34_17_n_9416 & mul_34_17_n_9287)));
 assign mul_34_17_n_9712 = ~(mul_34_17_n_11324 ^ mul_34_17_n_9454);
 assign mul_34_17_n_9711 = (mul_34_17_n_9221 ^ (mul_34_17_n_8768 ^ (mul_34_17_n_9223 ^ mul_34_17_n_9037)));
 assign mul_34_17_n_9710 = ((mul_34_17_n_9195 & mul_34_17_n_9295) | ((mul_34_17_n_9195 & mul_34_17_n_9351)
    | (mul_34_17_n_9351 & mul_34_17_n_9295)));
 assign mul_34_17_n_9709 = ((mul_34_17_n_11322 & mul_34_17_n_9427) | ((mul_34_17_n_11322 & mul_34_17_n_11318)
    | (mul_34_17_n_11318 & mul_34_17_n_9427)));
 assign mul_34_17_n_9706 = ~(mul_34_17_n_9508 ^ mul_34_17_n_9367);
 assign mul_34_17_n_9684 = ~mul_34_17_n_9683;
 assign mul_34_17_n_9681 = ~mul_34_17_n_9682;
 assign mul_34_17_n_9676 = ~mul_34_17_n_9675;
 assign mul_34_17_n_9672 = ~mul_34_17_n_11300;
 assign mul_34_17_n_9666 = ~mul_34_17_n_9667;
 assign mul_34_17_n_9658 = ~mul_34_17_n_9657;
 assign mul_34_17_n_9653 = ((mul_34_17_n_9190 & mul_34_17_n_285) | ((mul_34_17_n_9190 & mul_34_17_n_9191)
    | (mul_34_17_n_9191 & mul_34_17_n_285)));
 assign mul_34_17_n_9652 = ~(mul_34_17_n_9362 ^ mul_34_17_n_9438);
 assign mul_34_17_n_9651 = ~(mul_34_17_n_9083 | mul_34_17_n_356);
 assign mul_34_17_n_9650 = ~(mul_34_17_n_9510 & mul_34_17_n_9546);
 assign mul_34_17_n_9647 = ~(mul_34_17_n_357 | mul_34_17_n_9075);
 assign mul_34_17_n_9646 = ~((mul_34_17_n_9376 | mul_34_17_n_9304) & (mul_34_17_n_9087 | mul_34_17_n_8907));
 assign mul_34_17_n_9645 = ~(mul_34_17_n_9376 ^ mul_34_17_n_9304);
 assign mul_34_17_n_9644 = ~(mul_34_17_n_9526 & mul_34_17_n_9381);
 assign mul_34_17_n_9643 = ~(mul_34_17_n_9526 & mul_34_17_n_9305);
 assign mul_34_17_n_9641 = ~(mul_34_17_n_9523 & mul_34_17_n_9429);
 assign mul_34_17_n_9640 = ~(mul_34_17_n_9560 & mul_34_17_n_8953);
 assign mul_34_17_n_9639 = (mul_34_17_n_9225 ^ mul_34_17_n_9370);
 assign mul_34_17_n_9683 = ~(mul_34_17_n_9495 | mul_34_17_n_9211);
 assign mul_34_17_n_9638 = (mul_34_17_n_9115 ^ mul_34_17_n_9416);
 assign mul_34_17_n_9637 = ~(mul_34_17_n_279 ^ mul_34_17_n_9440);
 assign mul_34_17_n_9636 = ~(mul_34_17_n_9396 & (mul_34_17_n_9397 & (mul_34_17_n_9410 & mul_34_17_n_9308)));
 assign mul_34_17_n_9635 = (mul_34_17_n_9420 ^ mul_34_17_n_9424);
 assign mul_34_17_n_9634 = (mul_34_17_n_9220 ^ mul_34_17_n_9368);
 assign mul_34_17_n_9633 = ~(mul_34_17_n_9364 | mul_34_17_n_9501);
 assign mul_34_17_n_9632 = (mul_34_17_n_9228 ^ mul_34_17_n_277);
 assign mul_34_17_n_9682 = ((mul_34_17_n_9272 & mul_34_17_n_9360) | ((mul_34_17_n_9272 & mul_34_17_n_8849)
    | (mul_34_17_n_8849 & mul_34_17_n_9360)));
 assign mul_34_17_n_9631 = ~(mul_34_17_n_9535 & mul_34_17_n_9116);
 assign mul_34_17_n_9679 = ((mul_34_17_n_9171 & mul_34_17_n_9434) | ((mul_34_17_n_9171 & mul_34_17_n_9119)
    | (mul_34_17_n_9119 & mul_34_17_n_9434)));
 assign mul_34_17_n_9630 = ~(mul_34_17_n_9534 & mul_34_17_n_9117);
 assign mul_34_17_n_9678 = ((mul_34_17_n_272 & mul_34_17_n_9134) | ((mul_34_17_n_272 & mul_34_17_n_9216)
    | (mul_34_17_n_9216 & mul_34_17_n_9134)));
 assign mul_34_17_n_9677 = ((mul_34_17_n_9226 & mul_34_17_n_9230) | ((mul_34_17_n_9226 & mul_34_17_n_11328)
    | (mul_34_17_n_11328 & mul_34_17_n_9230)));
 assign mul_34_17_n_9675 = ~((mul_34_17_n_8879 | mul_34_17_n_8423) & (mul_34_17_n_9441 | mul_34_17_n_9131));
 assign mul_34_17_n_9629 = ~((mul_34_17_n_9444 & mul_34_17_n_9395) | (mul_34_17_n_9241 & mul_34_17_n_9069));
 assign mul_34_17_n_9674 = ((mul_34_17_n_9014 & mul_34_17_n_274) | ((mul_34_17_n_9014 & mul_34_17_n_8838)
    | (mul_34_17_n_8838 & mul_34_17_n_274)));
 assign mul_34_17_n_9670 = ~(mul_34_17_n_9479 & mul_34_17_n_9537);
 assign mul_34_17_n_9669 = ((mul_34_17_n_9267 & mul_34_17_n_11324) | ((mul_34_17_n_9267 & mul_34_17_n_9114)
    | (mul_34_17_n_9114 & mul_34_17_n_11324)));
 assign mul_34_17_n_9668 = ~(mul_34_17_n_9382 ^ mul_34_17_n_9269);
 assign mul_34_17_n_9667 = ~(mul_34_17_n_9192 ^ mul_34_17_n_9380);
 assign mul_34_17_n_9665 = ((mul_34_17_n_9178 & mul_34_17_n_8869) | ((mul_34_17_n_9178 & mul_34_17_n_8987)
    | (mul_34_17_n_8987 & mul_34_17_n_8869)));
 assign mul_34_17_n_9664 = ((mul_34_17_n_9269 & mul_34_17_n_9128) | ((mul_34_17_n_9269 & mul_34_17_n_8737)
    | (mul_34_17_n_8737 & mul_34_17_n_9128)));
 assign mul_34_17_n_9628 = (mul_34_17_n_9423 ^ mul_34_17_n_9296);
 assign mul_34_17_n_9663 = ((mul_34_17_n_9219 & mul_34_17_n_9367) | ((mul_34_17_n_9219 & mul_34_17_n_9045)
    | (mul_34_17_n_9045 & mul_34_17_n_9367)));
 assign mul_34_17_n_9662 = ((mul_34_17_n_268 & mul_34_17_n_9089) | ((mul_34_17_n_268 & mul_34_17_n_8984)
    | (mul_34_17_n_8984 & mul_34_17_n_9089)));
 assign mul_34_17_n_9661 = ~(mul_34_17_n_9289 ^ mul_34_17_n_9389);
 assign mul_34_17_n_9660 = ((mul_34_17_n_9275 & mul_34_17_n_8936) | ((mul_34_17_n_9275 & mul_34_17_n_9098)
    | (mul_34_17_n_9098 & mul_34_17_n_8936)));
 assign mul_34_17_n_9659 = ~((mul_34_17_n_9107 & (~mul_34_17_n_8925 & ~mul_34_17_n_9208)) | ((mul_34_17_n_9106
    & (mul_34_17_n_8925 & ~mul_34_17_n_9208)) | (mul_34_17_n_9401 & mul_34_17_n_9208)));
 assign mul_34_17_n_9657 = ~(mul_34_17_n_9383 ^ mul_34_17_n_8919);
 assign mul_34_17_n_9656 = ((mul_34_17_n_9215 & mul_34_17_n_9202) | ((mul_34_17_n_9215 & mul_34_17_n_9044)
    | (mul_34_17_n_9044 & mul_34_17_n_9202)));
 assign mul_34_17_n_9655 = ((mul_34_17_n_9192 & mul_34_17_n_11332) | ((mul_34_17_n_9192 & mul_34_17_n_9111)
    | (mul_34_17_n_9111 & mul_34_17_n_11332)));
 assign mul_34_17_n_9654 = ((mul_34_17_n_9163 & mul_34_17_n_9023) | ((mul_34_17_n_9163 & mul_34_17_n_8752)
    | (mul_34_17_n_8752 & mul_34_17_n_9023)));
 assign mul_34_17_n_9624 = ~mul_34_17_n_9625;
 assign mul_34_17_n_9623 = ~mul_34_17_n_9622;
 assign mul_34_17_n_9620 = ~mul_34_17_n_9621;
 assign mul_34_17_n_9612 = ~mul_34_17_n_11302;
 assign mul_34_17_n_9608 = ~mul_34_17_n_9607;
 assign mul_34_17_n_9605 = ~mul_34_17_n_9604;
 assign mul_34_17_n_9593 = ~mul_34_17_n_9592;
 assign mul_34_17_n_9589 = ~mul_34_17_n_9590;
 assign mul_34_17_n_9588 = ~mul_34_17_n_9587;
 assign mul_34_17_n_9580 = ~mul_34_17_n_9581;
 assign mul_34_17_n_9579 = ~(mul_34_17_n_9081 | mul_34_17_n_9521);
 assign mul_34_17_n_9578 = ~(mul_34_17_n_8880 ^ (mul_34_17_n_8385 ^ (mul_34_17_n_9043 ^ mul_34_17_n_8680)));
 assign mul_34_17_n_9572 = ((mul_34_17_n_9419 | mul_34_17_n_8998) & (mul_34_17_n_9170 | mul_34_17_n_8831));
 assign mul_34_17_n_9570 = ~(mul_34_17_n_9163 ^ mul_34_17_n_9345);
 assign mul_34_17_n_9569 = ~(mul_34_17_n_9188 ^ mul_34_17_n_9353);
 assign mul_34_17_n_9627 = ~(mul_34_17_n_9313 ^ mul_34_17_n_8942);
 assign mul_34_17_n_9626 = ~(mul_34_17_n_9193 ^ mul_34_17_n_280);
 assign mul_34_17_n_9625 = (mul_34_17_n_9427 ^ mul_34_17_n_11318);
 assign mul_34_17_n_9622 = ~(mul_34_17_n_9314 ^ mul_34_17_n_9147);
 assign mul_34_17_n_9568 = ~(mul_34_17_n_9333 ^ mul_34_17_n_9196);
 assign mul_34_17_n_9621 = (mul_34_17_n_9282 ^ mul_34_17_n_9349);
 assign mul_34_17_n_9567 = (mul_34_17_n_8849 ^ mul_34_17_n_9360);
 assign mul_34_17_n_9566 = (mul_34_17_n_290 ^ mul_34_17_n_9187);
 assign mul_34_17_n_9619 = ((mul_34_17_n_270 & mul_34_17_n_9262) | ((mul_34_17_n_270 & mul_34_17_n_8999)
    | (mul_34_17_n_8999 & mul_34_17_n_9262)));
 assign mul_34_17_n_9618 = ~(mul_34_17_n_9384 ^ mul_34_17_n_9123);
 assign mul_34_17_n_9617 = ~(mul_34_17_n_9345 ^ mul_34_17_n_9163);
 assign mul_34_17_n_9565 = ~(mul_34_17_n_9351 ^ mul_34_17_n_9195);
 assign mul_34_17_n_9616 = ~(mul_34_17_n_9035 ^ mul_34_17_n_9379);
 assign mul_34_17_n_9615 = ~(mul_34_17_n_9318 ^ mul_34_17_n_9090);
 assign mul_34_17_n_9564 = (mul_34_17_n_285 ^ mul_34_17_n_9190);
 assign mul_34_17_n_9614 = (mul_34_17_n_9415 ^ mul_34_17_n_9180);
 assign mul_34_17_n_9563 = (mul_34_17_n_9340 ^ mul_34_17_n_9301);
 assign mul_34_17_n_9562 = ~(mul_34_17_n_9316 ^ mul_34_17_n_8992);
 assign mul_34_17_n_9611 = ((mul_34_17_n_9173 & mul_34_17_n_9021) | ((mul_34_17_n_9173 & mul_34_17_n_9018)
    | (mul_34_17_n_9018 & mul_34_17_n_9021)));
 assign mul_34_17_n_9610 = ~(mul_34_17_n_9386 ^ mul_34_17_n_9277);
 assign mul_34_17_n_9609 = ((mul_34_17_n_9176 & mul_34_17_n_9205) | ((mul_34_17_n_9176 & mul_34_17_n_9004)
    | (mul_34_17_n_9004 & mul_34_17_n_9205)));
 assign mul_34_17_n_9607 = ((mul_34_17_n_9184 & mul_34_17_n_9285) | ((mul_34_17_n_9184 & mul_34_17_n_241)
    | (mul_34_17_n_241 & mul_34_17_n_9285)));
 assign mul_34_17_n_9606 = ((mul_34_17_n_9268 & mul_34_17_n_9260) | ((mul_34_17_n_9268 & mul_34_17_n_264)
    | (mul_34_17_n_264 & mul_34_17_n_9260)));
 assign mul_34_17_n_9604 = ~(mul_34_17_n_8985 ^ mul_34_17_n_9355);
 assign mul_34_17_n_9602 = ((mul_34_17_n_9186 & mul_34_17_n_9299) | ((mul_34_17_n_9186 & mul_34_17_n_9108)
    | (mul_34_17_n_9108 & mul_34_17_n_9299)));
 assign mul_34_17_n_9601 = ((mul_34_17_n_9169 & mul_34_17_n_9291) | ((mul_34_17_n_9169 & mul_34_17_n_9102)
    | (mul_34_17_n_9102 & mul_34_17_n_9291)));
 assign mul_34_17_n_9600 = ~(mul_34_17_n_9214 ^ mul_34_17_n_9320);
 assign mul_34_17_n_9599 = ((mul_34_17_n_9183 & mul_34_17_n_9027) | ((mul_34_17_n_9183 & mul_34_17_n_9013)
    | (mul_34_17_n_9013 & mul_34_17_n_9027)));
 assign mul_34_17_n_9598 = ~(mul_34_17_n_9275 ^ mul_34_17_n_9319);
 assign mul_34_17_n_9597 = ((mul_34_17_n_361 & mul_34_17_n_8553) | (mul_34_17_n_9404 & mul_34_17_n_8213));
 assign mul_34_17_n_9596 = ~(mul_34_17_n_9183 ^ mul_34_17_n_9312);
 assign mul_34_17_n_9595 = ((mul_34_17_n_9209 & mul_34_17_n_9263) | ((mul_34_17_n_9209 & mul_34_17_n_8829)
    | (mul_34_17_n_8829 & mul_34_17_n_9263)));
 assign mul_34_17_n_9594 = ~(mul_34_17_n_9315 ^ mul_34_17_n_9173);
 assign mul_34_17_n_9592 = (mul_34_17_n_9118 ^ mul_34_17_n_9373);
 assign mul_34_17_n_9591 = ((mul_34_17_n_9270 & mul_34_17_n_9292) | ((mul_34_17_n_9270 & mul_34_17_n_9093)
    | (mul_34_17_n_9093 & mul_34_17_n_9292)));
 assign mul_34_17_n_9590 = ((mul_34_17_n_9207 & mul_34_17_n_9261) | ((mul_34_17_n_9207 & mul_34_17_n_8982)
    | (mul_34_17_n_8982 & mul_34_17_n_9261)));
 assign mul_34_17_n_9587 = ((mul_34_17_n_260 & mul_34_17_n_9294) | ((mul_34_17_n_260 & mul_34_17_n_9001)
    | (mul_34_17_n_9001 & mul_34_17_n_9294)));
 assign mul_34_17_n_9585 = ~(mul_34_17_n_9206 ^ mul_34_17_n_9378);
 assign mul_34_17_n_9584 = ~((mul_34_17_n_8487 & (~mul_34_17_n_9113 & ~mul_34_17_n_9311)) | ((mul_34_17_n_8488
    & (mul_34_17_n_9113 & ~mul_34_17_n_9311)) | (mul_34_17_n_9433 & mul_34_17_n_9311)));
 assign mul_34_17_n_9583 = ((mul_34_17_n_9279 & mul_34_17_n_9288) | ((mul_34_17_n_9279 & mul_34_17_n_8927)
    | (mul_34_17_n_8927 & mul_34_17_n_9288)));
 assign mul_34_17_n_9582 = ~(mul_34_17_n_9317 ^ mul_34_17_n_9110);
 assign mul_34_17_n_9581 = (mul_34_17_n_9372 ^ mul_34_17_n_8618);
 assign mul_34_17_n_9552 = ~mul_34_17_n_9551;
 assign mul_34_17_n_9534 = ~mul_34_17_n_9535;
 assign mul_34_17_n_9525 = ~mul_34_17_n_9526;
 assign mul_34_17_n_9524 = ~(mul_34_17_n_0 ^ mul_34_17_n_8543);
 assign mul_34_17_n_9523 = ~(mul_34_17_n_9348 & mul_34_17_n_9281);
 assign mul_34_17_n_9522 = ~(mul_34_17_n_9349 & mul_34_17_n_9282);
 assign mul_34_17_n_9521 = (mul_34_17_n_9260 ^ mul_34_17_n_264);
 assign mul_34_17_n_9520 = ~(mul_34_17_n_358 | mul_34_17_n_8910);
 assign mul_34_17_n_9519 = ~(mul_34_17_n_9256 | mul_34_17_n_9407);
 assign mul_34_17_n_9518 = ~(mul_34_17_n_9226 ^ mul_34_17_n_11328);
 assign mul_34_17_n_9517 = ~(mul_34_17_n_8934 | (mul_34_17_n_9136 | (mul_34_17_n_9131 | mul_34_17_n_9132)));
 assign mul_34_17_n_9561 = ~(mul_34_17_n_9377 | mul_34_17_n_9231);
 assign mul_34_17_n_9515 = ((mul_34_17_n_8165 & mul_34_17_n_9302) | ((mul_34_17_n_8165 & mul_34_17_n_8070)
    | (mul_34_17_n_8070 & mul_34_17_n_9302)));
 assign mul_34_17_n_9560 = ((mul_34_17_n_8842 | mul_34_17_n_8912) & (mul_34_17_n_271 | mul_34_17_n_9105));
 assign mul_34_17_n_9514 = ~(mul_34_17_n_9387 | mul_34_17_n_8898);
 assign mul_34_17_n_9513 = (mul_34_17_n_9291 ^ mul_34_17_n_9102);
 assign mul_34_17_n_9559 = ~(mul_34_17_n_9266 ^ mul_34_17_n_8736);
 assign mul_34_17_n_9512 = ~(mul_34_17_n_272 ^ mul_34_17_n_9216);
 assign mul_34_17_n_9511 = ~(mul_34_17_n_9225 & mul_34_17_n_9370);
 assign mul_34_17_n_9558 = ((mul_34_17_n_9017 & mul_34_17_n_9031) | ((mul_34_17_n_9017 & mul_34_17_n_8993)
    | (mul_34_17_n_8993 & mul_34_17_n_9031)));
 assign mul_34_17_n_9557 = ~(mul_34_17_n_9288 ^ mul_34_17_n_9279);
 assign mul_34_17_n_9510 = ~(mul_34_17_n_9224 & mul_34_17_n_9371);
 assign mul_34_17_n_9556 = ((mul_34_17_n_8924 & mul_34_17_n_9208) | ((mul_34_17_n_8924 & mul_34_17_n_9107)
    | (mul_34_17_n_9107 & mul_34_17_n_9208)));
 assign mul_34_17_n_9509 = ((mul_34_17_n_8845 & mul_34_17_n_9298) | ((mul_34_17_n_8845 & mul_34_17_n_8619)
    | (mul_34_17_n_8619 & mul_34_17_n_9298)));
 assign mul_34_17_n_9555 = ((mul_34_17_n_362 & mul_34_17_n_9277) | ((mul_34_17_n_362 & mul_34_17_n_8732)
    | (mul_34_17_n_8732 & mul_34_17_n_9277)));
 assign mul_34_17_n_9508 = ~(mul_34_17_n_9219 ^ mul_34_17_n_9045);
 assign mul_34_17_n_9507 = ~(mul_34_17_n_9215 ^ mul_34_17_n_9044);
 assign mul_34_17_n_9554 = ((mul_34_17_n_9110 & mul_34_17_n_9030) | ((mul_34_17_n_9110 & mul_34_17_n_8644)
    | (mul_34_17_n_8644 & mul_34_17_n_9030)));
 assign mul_34_17_n_9553 = ~(mul_34_17_n_9293 ^ mul_34_17_n_8988);
 assign mul_34_17_n_9506 = ~(mul_34_17_n_9363 | mul_34_17_n_9437);
 assign mul_34_17_n_9505 = ~(mul_34_17_n_9140 ^ mul_34_17_n_8432);
 assign mul_34_17_n_9551 = ((mul_34_17_n_8989 & mul_34_17_n_9293) | ((mul_34_17_n_8989 & mul_34_17_n_9099)
    | (mul_34_17_n_9099 & mul_34_17_n_9293)));
 assign mul_34_17_n_9550 = ((mul_34_17_n_9112 & mul_34_17_n_9214) | ((mul_34_17_n_9112 & mul_34_17_n_8852)
    | (mul_34_17_n_8852 & mul_34_17_n_9214)));
 assign mul_34_17_n_9549 = ((mul_34_17_n_9101 & mul_34_17_n_9289) | ((mul_34_17_n_9101 & mul_34_17_n_8928)
    | (mul_34_17_n_8928 & mul_34_17_n_9289)));
 assign mul_34_17_n_9548 = ~((mul_34_17_n_8646 & (~mul_34_17_n_8840 & ~mul_34_17_n_9198)) | ((mul_34_17_n_8647
    & (mul_34_17_n_8840 & ~mul_34_17_n_9198)) | (mul_34_17_n_9243 & mul_34_17_n_9198)));
 assign mul_34_17_n_9547 = ((mul_34_17_n_8878 & mul_34_17_n_9206) | ((mul_34_17_n_8878 & mul_34_17_n_9040)
    | (mul_34_17_n_9040 & mul_34_17_n_9206)));
 assign mul_34_17_n_9546 = ((mul_34_17_n_11346 & mul_34_17_n_9200) | ((mul_34_17_n_11346 & mul_34_17_n_9104)
    | (mul_34_17_n_9104 & mul_34_17_n_9200)));
 assign mul_34_17_n_9545 = ((mul_34_17_n_9002 & mul_34_17_n_9046) | ((mul_34_17_n_9002 & mul_34_17_n_8645)
    | (mul_34_17_n_8645 & mul_34_17_n_9046)));
 assign mul_34_17_n_9544 = ~(mul_34_17_n_11619 ^ (mul_34_17_n_8745 ^ (mul_34_17_n_8570 ^ mul_34_17_n_8261)));
 assign mul_34_17_n_9543 = ~(mul_34_17_n_9363 & mul_34_17_n_9437);
 assign mul_34_17_n_9542 = ((mul_34_17_n_9039 & mul_34_17_n_9035) | ((mul_34_17_n_9039 & mul_34_17_n_9041)
    | (mul_34_17_n_9041 & mul_34_17_n_9035)));
 assign mul_34_17_n_9541 = ~(mul_34_17_n_267 ^ mul_34_17_n_9095);
 assign mul_34_17_n_9540 = ((mul_34_17_n_8839 & mul_34_17_n_9197) | ((mul_34_17_n_8839 & mul_34_17_n_8647)
    | (mul_34_17_n_8647 & mul_34_17_n_9197)));
 assign mul_34_17_n_9539 = ((mul_34_17_n_9109 & mul_34_17_n_11340) | ((mul_34_17_n_9109 & mul_34_17_n_9118)
    | (mul_34_17_n_9118 & mul_34_17_n_11340)));
 assign mul_34_17_n_9538 = ((mul_34_17_n_9038 & mul_34_17_n_9123) | ((mul_34_17_n_9038 & mul_34_17_n_263)
    | (mul_34_17_n_263 & mul_34_17_n_9123)));
 assign mul_34_17_n_9537 = ~((mul_34_17_n_8997 | mul_34_17_n_8244) & (mul_34_17_n_8942 | mul_34_17_n_9250));
 assign mul_34_17_n_9536 = ~(mul_34_17_n_9120 ^ mul_34_17_n_282);
 assign mul_34_17_n_9535 = ~(mul_34_17_n_9236 ^ mul_34_17_n_8539);
 assign mul_34_17_n_9533 = ((mul_34_17_n_9090 & mul_34_17_n_9028) | ((mul_34_17_n_9090 & mul_34_17_n_257)
    | (mul_34_17_n_257 & mul_34_17_n_9028)));
 assign mul_34_17_n_9532 = ((mul_34_17_n_9122 & mul_34_17_n_9210) | ((mul_34_17_n_9122 & mul_34_17_n_9019)
    | (mul_34_17_n_9019 & mul_34_17_n_9210)));
 assign mul_34_17_n_9531 = ((mul_34_17_n_9003 & mul_34_17_n_9025) | ((mul_34_17_n_9003 & mul_34_17_n_8985)
    | (mul_34_17_n_8985 & mul_34_17_n_9025)));
 assign mul_34_17_n_9530 = ~((mul_34_17_n_9080 & mul_34_17_n_8803) | (mul_34_17_n_9252 & mul_34_17_n_8477));
 assign mul_34_17_n_9529 = ~(mul_34_17_n_9233 ^ mul_34_17_n_8758);
 assign mul_34_17_n_9528 = ~(mul_34_17_n_9234 ^ mul_34_17_n_8692);
 assign mul_34_17_n_9527 = ((mul_34_17_n_9086 | mul_34_17_n_269) & (mul_34_17_n_9255 | mul_34_17_n_8717));
 assign mul_34_17_n_9526 = ~(mul_34_17_n_9071 & (mul_34_17_n_8950 & (mul_34_17_n_9248 & mul_34_17_n_9251)));
 assign mul_34_17_n_9494 = ~mul_34_17_n_9495;
 assign mul_34_17_n_9478 = ~mul_34_17_n_9477;
 assign mul_34_17_n_9461 = ~(mul_34_17_n_9185 ^ mul_34_17_n_8827);
 assign mul_34_17_n_9460 = (mul_34_17_n_264 ^ mul_34_17_n_9260);
 assign mul_34_17_n_9458 = ~(mul_34_17_n_9164 ^ mul_34_17_n_8602);
 assign mul_34_17_n_9457 = ~(mul_34_17_n_9284 ^ mul_34_17_n_266);
 assign mul_34_17_n_9456 = ((mul_34_17_n_8659 & mul_34_17_n_9203) | ((mul_34_17_n_8659 & mul_34_17_n_8373)
    | (mul_34_17_n_8373 & mul_34_17_n_9203)));
 assign mul_34_17_n_9455 = ~(mul_34_17_n_230 ^ (mul_34_17_n_8382 ^ (mul_34_17_n_8690 ^ mul_34_17_n_8511)));
 assign mul_34_17_n_9504 = (mul_34_17_n_9186 ^ mul_34_17_n_9108);
 assign mul_34_17_n_9454 = (mul_34_17_n_9267 ^ mul_34_17_n_9114);
 assign mul_34_17_n_9503 = ~(mul_34_17_n_265 ^ mul_34_17_n_8361);
 assign mul_34_17_n_9453 = (mul_34_17_n_9176 ^ mul_34_17_n_9004);
 assign mul_34_17_n_9502 = ~(mul_34_17_n_9105 ^ mul_34_17_n_271);
 assign mul_34_17_n_9501 = ~(mul_34_17_n_9185 ^ mul_34_17_n_8826);
 assign mul_34_17_n_9452 = (mul_34_17_n_9294 ^ mul_34_17_n_260);
 assign mul_34_17_n_9500 = ~(mul_34_17_n_9143 ^ mul_34_17_n_8741);
 assign mul_34_17_n_9451 = (mul_34_17_n_9270 ^ mul_34_17_n_9292);
 assign mul_34_17_n_9499 = ~(mul_34_17_n_9203 ^ mul_34_17_n_9138);
 assign mul_34_17_n_9498 = (mul_34_17_n_9178 ^ mul_34_17_n_8869);
 assign mul_34_17_n_9450 = ~(mul_34_17_n_9171 ^ mul_34_17_n_9119);
 assign mul_34_17_n_9449 = ~(mul_34_17_n_9285 ^ mul_34_17_n_241);
 assign mul_34_17_n_9448 = (mul_34_17_n_9210 ^ mul_34_17_n_9019);
 assign mul_34_17_n_9497 = ~(mul_34_17_n_9144 ^ mul_34_17_n_8931);
 assign mul_34_17_n_9495 = ~(mul_34_17_n_9148 ^ mul_34_17_n_8522);
 assign mul_34_17_n_9493 = ~(mul_34_17_n_9149 ^ mul_34_17_n_8854);
 assign mul_34_17_n_9447 = (mul_34_17_n_9221 ^ mul_34_17_n_8768);
 assign mul_34_17_n_9492 = ~(mul_34_17_n_9194 ^ mul_34_17_n_8597);
 assign mul_34_17_n_9491 = ~(mul_34_17_n_9151 ^ mul_34_17_n_9026);
 assign mul_34_17_n_9490 = ~(mul_34_17_n_9152 ^ mul_34_17_n_9011);
 assign mul_34_17_n_9489 = ~((mul_34_17_n_8761 & (~mul_34_17_n_8932 & ~mul_34_17_n_9127)) | ((mul_34_17_n_8760
    & (mul_34_17_n_8932 & ~mul_34_17_n_9127)) | (mul_34_17_n_9242 & mul_34_17_n_9127)));
 assign mul_34_17_n_9487 = ~(mul_34_17_n_9142 ^ mul_34_17_n_8846);
 assign mul_34_17_n_9485 = ~(mul_34_17_n_8738 ^ mul_34_17_n_9141);
 assign mul_34_17_n_9446 = ~(mul_34_17_n_9229 ^ mul_34_17_n_9297);
 assign mul_34_17_n_9483 = ~((mul_34_17_n_8721 & (~mul_34_17_n_8915 & ~mul_34_17_n_254)) | ((mul_34_17_n_8722
    & (mul_34_17_n_8915 & ~mul_34_17_n_254)) | (mul_34_17_n_9244 & mul_34_17_n_254)));
 assign mul_34_17_n_9482 = ~(mul_34_17_n_9150 ^ mul_34_17_n_9029);
 assign mul_34_17_n_9481 = ((mul_34_17_n_8991 & mul_34_17_n_11330) | ((mul_34_17_n_8991 & mul_34_17_n_8995)
    | (mul_34_17_n_8995 & mul_34_17_n_11330)));
 assign mul_34_17_n_9480 = ((mul_34_17_n_9091 & mul_34_17_n_11338) | ((mul_34_17_n_9091 & mul_34_17_n_8926)
    | (mul_34_17_n_8926 & mul_34_17_n_11338)));
 assign mul_34_17_n_9445 = ~(mul_34_17_n_9217 ^ mul_34_17_n_8859);
 assign mul_34_17_n_9479 = ~(mul_34_17_n_9218 ^ mul_34_17_n_8940);
 assign mul_34_17_n_9477 = ~(mul_34_17_n_9167 ^ mul_34_17_n_9174);
 assign mul_34_17_n_9476 = ~(mul_34_17_n_9146 ^ mul_34_17_n_9009);
 assign mul_34_17_n_9475 = ((mul_34_17_n_9007 & mul_34_17_n_11348) | ((mul_34_17_n_9007 & mul_34_17_n_8730)
    | (mul_34_17_n_8730 & mul_34_17_n_11348)));
 assign mul_34_17_n_9474 = (mul_34_17_n_270 ^ mul_34_17_n_8999);
 assign mul_34_17_n_9473 = ((mul_34_17_n_9011 & mul_34_17_n_11621) | ((mul_34_17_n_9011 & mul_34_17_n_8841)
    | (mul_34_17_n_8841 & mul_34_17_n_11621)));
 assign mul_34_17_n_9472 = ((mul_34_17_n_9088 & mul_34_17_n_267) | ((mul_34_17_n_9088 & mul_34_17_n_9096)
    | (mul_34_17_n_9096 & mul_34_17_n_267)));
 assign mul_34_17_n_9470 = ((mul_34_17_n_359 & mul_34_17_n_8801) | (mul_34_17_n_9240 & mul_34_17_n_8460));
 assign mul_34_17_n_9469 = ~(mul_34_17_n_9145 ^ mul_34_17_n_8254);
 assign mul_34_17_n_9468 = ((mul_34_17_n_9010 & mul_34_17_n_8874) | ((mul_34_17_n_9010 & mul_34_17_n_8633)
    | (mul_34_17_n_8633 & mul_34_17_n_8874)));
 assign mul_34_17_n_9467 = ~((mul_34_17_n_8601 & mul_34_17_n_8637) | (mul_34_17_n_9164 & mul_34_17_n_8909));
 assign mul_34_17_n_9466 = ~((mul_34_17_n_8595 & (~mul_34_17_n_8835 & ~mul_34_17_n_8662)) | ((mul_34_17_n_8594
    & (mul_34_17_n_8835 & ~mul_34_17_n_8662)) | (mul_34_17_n_9154 & mul_34_17_n_8662)));
 assign mul_34_17_n_9464 = ((mul_34_17_n_360 & mul_34_17_n_8670) | (mul_34_17_n_9245 & mul_34_17_n_8462));
 assign mul_34_17_n_9463 = ~(mul_34_17_n_9307 ^ mul_34_17_n_9092);
 assign mul_34_17_n_9462 = ~(mul_34_17_n_9238 ^ mul_34_17_n_8507);
 assign mul_34_17_n_9444 = ~mul_34_17_n_9394;
 assign mul_34_17_n_9437 = ~mul_34_17_n_9438;
 assign mul_34_17_n_9436 = ~mul_34_17_n_9435;
 assign mul_34_17_n_9431 = ~mul_34_17_n_9430;
 assign mul_34_17_n_9428 = ~mul_34_17_n_9429;
 assign mul_34_17_n_9421 = ~mul_34_17_n_9422;
 assign mul_34_17_n_9417 = ~mul_34_17_n_9418;
 assign mul_34_17_n_9410 = ((mul_34_17_n_8997 & mul_34_17_n_8244) | (mul_34_17_n_8709 & mul_34_17_n_8698));
 assign mul_34_17_n_9409 = ~(mul_34_17_n_9208 & mul_34_17_n_9237);
 assign mul_34_17_n_9407 = (mul_34_17_n_8986 ^ mul_34_17_n_8913);
 assign mul_34_17_n_9406 = ~(mul_34_17_n_9266 & mul_34_17_n_8736);
 assign mul_34_17_n_9405 = ~(mul_34_17_n_9266 | mul_34_17_n_8736);
 assign mul_34_17_n_9404 = ~(mul_34_17_n_361 | mul_34_17_n_8212);
 assign mul_34_17_n_9403 = ~(mul_34_17_n_236 ^ mul_34_17_n_8791);
 assign mul_34_17_n_9402 = (mul_34_17_n_8913 ^ mul_34_17_n_8986);
 assign mul_34_17_n_9401 = ~(mul_34_17_n_8925 ^ mul_34_17_n_9107);
 assign mul_34_17_n_9399 = ~(mul_34_17_n_9194 & mul_34_17_n_8597);
 assign mul_34_17_n_9398 = ~(mul_34_17_n_9194 | mul_34_17_n_8597);
 assign mul_34_17_n_9397 = ~(mul_34_17_n_9218 & mul_34_17_n_8940);
 assign mul_34_17_n_9396 = ~(mul_34_17_n_9076 & (mul_34_17_n_9077 & (mul_34_17_n_8708 & mul_34_17_n_8177)));
 assign mul_34_17_n_9395 = ~(mul_34_17_n_9203 & mul_34_17_n_9138);
 assign mul_34_17_n_9394 = ~(mul_34_17_n_9203 | mul_34_17_n_9138);
 assign mul_34_17_n_9393 = ~(mul_34_17_n_9170 & mul_34_17_n_8831);
 assign mul_34_17_n_9392 = ((mul_34_17_n_8845 & mul_34_17_n_8974) | ((mul_34_17_n_8845 & mul_34_17_n_8619)
    | (mul_34_17_n_8619 & mul_34_17_n_8974)));
 assign mul_34_17_n_9391 = ~(mul_34_17_n_271 & mul_34_17_n_9105);
 assign mul_34_17_n_9443 = ~(mul_34_17_n_9276 & mul_34_17_n_8914);
 assign mul_34_17_n_9390 = ~(mul_34_17_n_9276 | mul_34_17_n_8914);
 assign mul_34_17_n_9389 = (mul_34_17_n_8928 ^ mul_34_17_n_9101);
 assign mul_34_17_n_9387 = ~(mul_34_17_n_9275 | mul_34_17_n_9098);
 assign mul_34_17_n_9386 = (mul_34_17_n_362 ^ mul_34_17_n_8732);
 assign mul_34_17_n_9385 = ~(mul_34_17_n_9275 & mul_34_17_n_9098);
 assign mul_34_17_n_9384 = (mul_34_17_n_9038 ^ mul_34_17_n_263);
 assign mul_34_17_n_9383 = ~(mul_34_17_n_9125 ^ mul_34_17_n_8764);
 assign mul_34_17_n_9441 = ((mul_34_17_n_8688 | mul_34_17_n_8428) & (mul_34_17_n_8934 | mul_34_17_n_9065));
 assign mul_34_17_n_9382 = (mul_34_17_n_8737 ^ mul_34_17_n_9128);
 assign mul_34_17_n_9381 = ~(mul_34_17_n_9306 | mul_34_17_n_9131);
 assign mul_34_17_n_9380 = ~(mul_34_17_n_11332 ^ mul_34_17_n_9111);
 assign mul_34_17_n_9379 = (mul_34_17_n_9039 ^ mul_34_17_n_9041);
 assign mul_34_17_n_9378 = ~(mul_34_17_n_8878 ^ mul_34_17_n_9040);
 assign mul_34_17_n_9440 = ((mul_34_17_n_8914 & mul_34_17_n_11619) | ((mul_34_17_n_8914 & mul_34_17_n_8745)
    | (mul_34_17_n_8745 & mul_34_17_n_11619)));
 assign mul_34_17_n_9439 = ((mul_34_17_n_8931 & mul_34_17_n_8876) | ((mul_34_17_n_8931 & mul_34_17_n_8381)
    | (mul_34_17_n_8381 & mul_34_17_n_8876)));
 assign mul_34_17_n_9438 = ((mul_34_17_n_8865 & mul_34_17_n_8150) | ((mul_34_17_n_8865 & mul_34_17_n_8740)
    | (mul_34_17_n_8740 & mul_34_17_n_8150)));
 assign mul_34_17_n_9435 = ~(mul_34_17_n_8568 ^ (mul_34_17_n_8750 ^ (mul_34_17_n_8273 ^ mul_34_17_n_7739)));
 assign mul_34_17_n_9434 = ~((mul_34_17_n_8352 & (~mul_34_17_n_8655 & ~mul_34_17_n_275)) | ((mul_34_17_n_8353
    & (mul_34_17_n_8655 & ~mul_34_17_n_275)) | (mul_34_17_n_9066 & mul_34_17_n_275)));
 assign mul_34_17_n_9433 = ~(mul_34_17_n_9113 ^ mul_34_17_n_8487);
 assign mul_34_17_n_9377 = ~(mul_34_17_n_9226 | mul_34_17_n_11328);
 assign mul_34_17_n_9430 = ~(mul_34_17_n_9055 ^ mul_34_17_n_9124);
 assign mul_34_17_n_9429 = ~(mul_34_17_n_9053 ^ mul_34_17_n_8864);
 assign mul_34_17_n_9427 = ((mul_34_17_n_8894 & mul_34_17_n_8735) | ((mul_34_17_n_8894 & mul_34_17_n_8890)
    | (mul_34_17_n_8890 & mul_34_17_n_8735)));
 assign mul_34_17_n_9426 = ((mul_34_17_n_8920 & mul_34_17_n_9125) | ((mul_34_17_n_8920 & mul_34_17_n_8765)
    | (mul_34_17_n_8765 & mul_34_17_n_9125)));
 assign mul_34_17_n_9425 = ((mul_34_17_n_8802 & mul_34_17_n_9129) | ((mul_34_17_n_8802 & mul_34_17_n_11350)
    | (mul_34_17_n_11350 & mul_34_17_n_9129)));
 assign mul_34_17_n_9424 = ((mul_34_17_n_8761 & mul_34_17_n_9126) | ((mul_34_17_n_8761 & mul_34_17_n_8932)
    | (mul_34_17_n_8932 & mul_34_17_n_9126)));
 assign mul_34_17_n_9423 = ~(mul_34_17_n_9049 ^ mul_34_17_n_8549);
 assign mul_34_17_n_9422 = ((mul_34_17_n_273 & mul_34_17_n_8834) | ((mul_34_17_n_273 & mul_34_17_n_8724)
    | (mul_34_17_n_8724 & mul_34_17_n_8834)));
 assign mul_34_17_n_9420 = ~(mul_34_17_n_9050 ^ mul_34_17_n_8943);
 assign mul_34_17_n_9419 = ((mul_34_17_n_8656 & mul_34_17_n_9034) | ((mul_34_17_n_8656 & mul_34_17_n_8353)
    | (mul_34_17_n_8353 & mul_34_17_n_9034)));
 assign mul_34_17_n_9418 = ((mul_34_17_n_8923 & mul_34_17_n_11342) | ((mul_34_17_n_8923 & mul_34_17_n_8640)
    | (mul_34_17_n_8640 & mul_34_17_n_11342)));
 assign mul_34_17_n_9416 = ~(mul_34_17_n_9054 ^ mul_34_17_n_8512);
 assign mul_34_17_n_9415 = ~((mul_34_17_n_8628 & (~mul_34_17_n_8626 & ~mul_34_17_n_8872)) | ((mul_34_17_n_8627
    & (mul_34_17_n_8626 & ~mul_34_17_n_8872)) | (mul_34_17_n_8975 & mul_34_17_n_8872)));
 assign mul_34_17_n_9411 = ((mul_34_17_n_8930 & mul_34_17_n_8949) | ((mul_34_17_n_8930 & mul_34_17_n_8738)
    | (mul_34_17_n_8738 & mul_34_17_n_8949)));
 assign mul_34_17_n_9371 = ~mul_34_17_n_9370;
 assign mul_34_17_n_9365 = ~mul_34_17_n_9364;
 assign mul_34_17_n_9362 = ~mul_34_17_n_9363;
 assign mul_34_17_n_9357 = ~mul_34_17_n_11322;
 assign mul_34_17_n_9349 = ~mul_34_17_n_9348;
 assign mul_34_17_n_9347 = ~mul_34_17_n_9346;
 assign mul_34_17_n_9339 = ~mul_34_17_n_9338;
 assign mul_34_17_n_9325 = ~mul_34_17_n_278;
 assign mul_34_17_n_9320 = (mul_34_17_n_9112 ^ mul_34_17_n_8852);
 assign mul_34_17_n_9376 = ~((mul_34_17_n_8396 & (~mul_34_17_n_7681 & ~mul_34_17_n_8956)) | ((mul_34_17_n_8397
    & (mul_34_17_n_7681 & ~mul_34_17_n_8956)) | (mul_34_17_n_8865 & mul_34_17_n_8956)));
 assign mul_34_17_n_9319 = (mul_34_17_n_9098 ^ mul_34_17_n_8936);
 assign mul_34_17_n_9375 = ((mul_34_17_n_8827 & mul_34_17_n_11344) | ((mul_34_17_n_8827 & mul_34_17_n_8631)
    | (mul_34_17_n_8631 & mul_34_17_n_11344)));
 assign mul_34_17_n_9318 = (mul_34_17_n_9028 ^ mul_34_17_n_257);
 assign mul_34_17_n_9317 = (mul_34_17_n_9030 ^ mul_34_17_n_8644);
 assign mul_34_17_n_9316 = (mul_34_17_n_8492 ^ mul_34_17_n_9006);
 assign mul_34_17_n_9374 = ((mul_34_17_n_259 & mul_34_17_n_8940) | ((mul_34_17_n_259 & mul_34_17_n_256)
    | (mul_34_17_n_256 & mul_34_17_n_8940)));
 assign mul_34_17_n_9373 = ~(mul_34_17_n_11340 ^ mul_34_17_n_9109);
 assign mul_34_17_n_9372 = ~(mul_34_17_n_9033 ^ mul_34_17_n_11364);
 assign mul_34_17_n_9315 = ~(mul_34_17_n_9021 ^ mul_34_17_n_9018);
 assign mul_34_17_n_9314 = (mul_34_17_n_9005 ^ mul_34_17_n_8851);
 assign mul_34_17_n_9370 = ~(mul_34_17_n_8971 ^ mul_34_17_n_8379);
 assign mul_34_17_n_9369 = ((mul_34_17_n_8621 & mul_34_17_n_9024) | ((mul_34_17_n_8621 & mul_34_17_n_8247)
    | (mul_34_17_n_8247 & mul_34_17_n_9024)));
 assign mul_34_17_n_9368 = ~(mul_34_17_n_8954 ^ mul_34_17_n_8657);
 assign mul_34_17_n_9313 = ~(mul_34_17_n_8997 ^ mul_34_17_n_8244);
 assign mul_34_17_n_9312 = ~(mul_34_17_n_9013 ^ mul_34_17_n_9027);
 assign mul_34_17_n_9311 = ~(mul_34_17_n_9130 ^ mul_34_17_n_8929);
 assign mul_34_17_n_9310 = (mul_34_17_n_11330 ^ mul_34_17_n_8991);
 assign mul_34_17_n_9367 = ((mul_34_17_n_240 & mul_34_17_n_8779) | ((mul_34_17_n_240 & mul_34_17_n_8508)
    | (mul_34_17_n_8508 & mul_34_17_n_8779)));
 assign mul_34_17_n_9366 = ~((mul_34_17_n_8719 & (~mul_34_17_n_8600 & ~mul_34_17_n_8948)) | ((mul_34_17_n_8720
    & (mul_34_17_n_8600 & ~mul_34_17_n_8948)) | (mul_34_17_n_9068 & mul_34_17_n_8948)));
 assign mul_34_17_n_9364 = ~(mul_34_17_n_8969 ^ mul_34_17_n_8638);
 assign mul_34_17_n_9363 = ~(mul_34_17_n_9024 ^ mul_34_17_n_8960);
 assign mul_34_17_n_9361 = ~(mul_34_17_n_9012 ^ mul_34_17_n_8917);
 assign mul_34_17_n_9360 = ~(mul_34_17_n_8957 ^ mul_34_17_n_8939);
 assign mul_34_17_n_9359 = ((mul_34_17_n_8762 & mul_34_17_n_9124) | ((mul_34_17_n_8762 & mul_34_17_n_8763)
    | (mul_34_17_n_8763 & mul_34_17_n_9124)));
 assign mul_34_17_n_9356 = ((mul_34_17_n_8922 & mul_34_17_n_8609) | ((mul_34_17_n_8922 & mul_34_17_n_8723)
    | (mul_34_17_n_8723 & mul_34_17_n_8609)));
 assign mul_34_17_n_9309 = (mul_34_17_n_9042 ^ mul_34_17_n_8375);
 assign mul_34_17_n_9355 = (mul_34_17_n_9025 ^ mul_34_17_n_9003);
 assign mul_34_17_n_9354 = ((mul_34_17_n_8854 & mul_34_17_n_8805) | ((mul_34_17_n_8854 & mul_34_17_n_8575)
    | (mul_34_17_n_8575 & mul_34_17_n_8805)));
 assign mul_34_17_n_9353 = ~(mul_34_17_n_8962 ^ mul_34_17_n_8406);
 assign mul_34_17_n_9352 = ~(mul_34_17_n_8955 ^ mul_34_17_n_8370);
 assign mul_34_17_n_9351 = ~(mul_34_17_n_8958 ^ mul_34_17_n_8684);
 assign mul_34_17_n_9350 = ~(mul_34_17_n_8964 ^ mul_34_17_n_8789);
 assign mul_34_17_n_9348 = ~(mul_34_17_n_9056 ^ mul_34_17_n_8500);
 assign mul_34_17_n_9346 = ~(mul_34_17_n_8965 ^ mul_34_17_n_8363);
 assign mul_34_17_n_9345 = ~(mul_34_17_n_9023 ^ mul_34_17_n_8752);
 assign mul_34_17_n_9344 = ((mul_34_17_n_8635 & mul_34_17_n_9033) | ((mul_34_17_n_8635 & mul_34_17_n_8618)
    | (mul_34_17_n_8618 & mul_34_17_n_9033)));
 assign mul_34_17_n_9343 = ~(mul_34_17_n_9052 ^ mul_34_17_n_8393);
 assign mul_34_17_n_9342 = (mul_34_17_n_9043 ^ mul_34_17_n_8680);
 assign mul_34_17_n_9341 = ~(mul_34_17_n_8591 ^ (mul_34_17_n_8603 ^ (mul_34_17_n_8426 ^ mul_34_17_n_7535)));
 assign mul_34_17_n_9340 = ~(mul_34_17_n_8970 ^ mul_34_17_n_8232);
 assign mul_34_17_n_9338 = ((mul_34_17_n_230 & mul_34_17_n_8830) | ((mul_34_17_n_230 & mul_34_17_n_8382)
    | (mul_34_17_n_8382 & mul_34_17_n_8830)));
 assign mul_34_17_n_9337 = ((mul_34_17_n_244 & mul_34_17_n_9029) | ((mul_34_17_n_244 & mul_34_17_n_8625)
    | (mul_34_17_n_8625 & mul_34_17_n_9029)));
 assign mul_34_17_n_9336 = ~(mul_34_17_n_9048 ^ mul_34_17_n_8359);
 assign mul_34_17_n_9334 = ((mul_34_17_n_8933 & mul_34_17_n_8866) | ((mul_34_17_n_8933 & mul_34_17_n_8847)
    | (mul_34_17_n_8847 & mul_34_17_n_8866)));
 assign mul_34_17_n_9333 = ~(mul_34_17_n_9057 ^ mul_34_17_n_8529);
 assign mul_34_17_n_9332 = ~(mul_34_17_n_8959 ^ mul_34_17_n_8369);
 assign mul_34_17_n_9331 = ~((mul_34_17_n_11368 & (~mul_34_17_n_8734 & ~mul_34_17_n_8746)) | ((mul_34_17_n_8605
    & (mul_34_17_n_8734 & ~mul_34_17_n_8746)) | (mul_34_17_n_8981 & mul_34_17_n_8746)));
 assign mul_34_17_n_9330 = ((mul_34_17_n_8853 & mul_34_17_n_9026) | ((mul_34_17_n_8853 & mul_34_17_n_8650)
    | (mul_34_17_n_8650 & mul_34_17_n_9026)));
 assign mul_34_17_n_9329 = ((mul_34_17_n_8843 & mul_34_17_n_8867) | ((mul_34_17_n_8843 & mul_34_17_n_8596)
    | (mul_34_17_n_8596 & mul_34_17_n_8867)));
 assign mul_34_17_n_9328 = ~(mul_34_17_n_8961 ^ mul_34_17_n_8877);
 assign mul_34_17_n_9327 = ((mul_34_17_n_254 & mul_34_17_n_8915) | ((mul_34_17_n_254 & mul_34_17_n_8721)
    | (mul_34_17_n_8721 & mul_34_17_n_8915)));
 assign mul_34_17_n_9326 = ~(mul_34_17_n_9051 ^ mul_34_17_n_8677);
 assign mul_34_17_n_9308 = ~mul_34_17_n_9258;
 assign mul_34_17_n_9306 = ~mul_34_17_n_9305;
 assign mul_34_17_n_9300 = ~mul_34_17_n_9299;
 assign mul_34_17_n_9298 = ~mul_34_17_n_9297;
 assign mul_34_17_n_9282 = ~mul_34_17_n_9281;
 assign mul_34_17_n_9259 = ~(mul_34_17_n_8879 ^ mul_34_17_n_8423);
 assign mul_34_17_n_9258 = ~(mul_34_17_n_8997 | mul_34_17_n_8244);
 assign mul_34_17_n_9257 = ~(mul_34_17_n_9097 & mul_34_17_n_8727);
 assign mul_34_17_n_9256 = ~(mul_34_17_n_9097 | mul_34_17_n_8727);
 assign mul_34_17_n_9255 = ~(mul_34_17_n_9067 & mul_34_17_n_8716);
 assign mul_34_17_n_9254 = ~(mul_34_17_n_9012 | mul_34_17_n_8917);
 assign mul_34_17_n_9253 = ~(mul_34_17_n_9012 & mul_34_17_n_8917);
 assign mul_34_17_n_9252 = ~(mul_34_17_n_8976 | mul_34_17_n_8476);
 assign mul_34_17_n_9251 = ~(mul_34_17_n_8799 & (mul_34_17_n_8280 & (mul_34_17_n_8272 & mul_34_17_n_9137)));
 assign mul_34_17_n_9250 = ~(mul_34_17_n_8996 | mul_34_17_n_8243);
 assign mul_34_17_n_9249 = ~(mul_34_17_n_11334 ^ mul_34_17_n_8804);
 assign mul_34_17_n_9248 = ~(mul_34_17_n_9137 & mul_34_17_n_8792);
 assign mul_34_17_n_9245 = ~(mul_34_17_n_360 | mul_34_17_n_8463);
 assign mul_34_17_n_9244 = ~(mul_34_17_n_8571 ^ (mul_34_17_n_7745 ^ (mul_34_17_n_8278 ^ mul_34_17_n_7566)));
 assign mul_34_17_n_9243 = ~(mul_34_17_n_8427 ^ (mul_34_17_n_7858 ^ (mul_34_17_n_7066 ^ mul_34_17_n_8171)));
 assign mul_34_17_n_9242 = ~(mul_34_17_n_8275 ^ (mul_34_17_n_7767 ^ (mul_34_17_n_253 ^ mul_34_17_n_7734)));
 assign mul_34_17_n_9241 = ~(mul_34_17_n_9139 & mul_34_17_n_8940);
 assign mul_34_17_n_9240 = ~(mul_34_17_n_359 | mul_34_17_n_8461);
 assign mul_34_17_n_9239 = ((mul_34_17_n_8608 & mul_34_17_n_8448) | ((mul_34_17_n_8608 & mul_34_17_n_8331)
    | (mul_34_17_n_8331 & mul_34_17_n_8448)));
 assign mul_34_17_n_9307 = (mul_34_17_n_11338 ^ mul_34_17_n_8926);
 assign mul_34_17_n_9238 = (mul_34_17_n_8779 ^ mul_34_17_n_240);
 assign mul_34_17_n_9237 = ~(mul_34_17_n_8925 & mul_34_17_n_9106);
 assign mul_34_17_n_9236 = ~(mul_34_17_n_8941 ^ mul_34_17_n_8517);
 assign mul_34_17_n_9305 = ~(mul_34_17_n_8934 | mul_34_17_n_9136);
 assign mul_34_17_n_9235 = ~(mul_34_17_n_8924 & mul_34_17_n_9107);
 assign mul_34_17_n_9234 = ((mul_34_17_n_8728 & mul_34_17_n_8568) | ((mul_34_17_n_8728 & mul_34_17_n_8750)
    | (mul_34_17_n_8750 & mul_34_17_n_8568)));
 assign mul_34_17_n_9233 = ~(mul_34_17_n_8944 ^ mul_34_17_n_8759);
 assign mul_34_17_n_9304 = ((mul_34_17_n_8522 & mul_34_17_n_8873) | ((mul_34_17_n_8522 & mul_34_17_n_8248)
    | (mul_34_17_n_8248 & mul_34_17_n_8873)));
 assign mul_34_17_n_9303 = ((mul_34_17_n_8626 & mul_34_17_n_8872) | ((mul_34_17_n_8626 & mul_34_17_n_8628)
    | (mul_34_17_n_8628 & mul_34_17_n_8872)));
 assign mul_34_17_n_9302 = ~(mul_34_17_n_9062 & mul_34_17_n_8793);
 assign mul_34_17_n_9301 = ((mul_34_17_n_363 & mul_34_17_n_7945) | (mul_34_17_n_8903 & mul_34_17_n_7612));
 assign mul_34_17_n_9299 = ((mul_34_17_n_8742 & mul_34_17_n_11336) | ((mul_34_17_n_8742 & mul_34_17_n_8632)
    | (mul_34_17_n_8632 & mul_34_17_n_11336)));
 assign mul_34_17_n_9297 = ((mul_34_17_n_8610 & mul_34_17_n_8489) | ((mul_34_17_n_8610 & mul_34_17_n_7980)
    | (mul_34_17_n_7980 & mul_34_17_n_8489)));
 assign mul_34_17_n_9296 = ((mul_34_17_n_8753 & mul_34_17_n_11362) | ((mul_34_17_n_8753 & mul_34_17_n_8751)
    | (mul_34_17_n_8751 & mul_34_17_n_11362)));
 assign mul_34_17_n_9295 = ((mul_34_17_n_8687 & mul_34_17_n_8678) | ((mul_34_17_n_8687 & mul_34_17_n_8425)
    | (mul_34_17_n_8425 & mul_34_17_n_8678)));
 assign mul_34_17_n_9294 = ((mul_34_17_n_8739 & mul_34_17_n_8773) | ((mul_34_17_n_8739 & mul_34_17_n_8140)
    | (mul_34_17_n_8140 & mul_34_17_n_8773)));
 assign mul_34_17_n_9293 = ~(mul_34_17_n_8887 ^ mul_34_17_n_8775);
 assign mul_34_17_n_9292 = ((mul_34_17_n_8733 & mul_34_17_n_8801) | ((mul_34_17_n_8733 & mul_34_17_n_8493)
    | (mul_34_17_n_8493 & mul_34_17_n_8801)));
 assign mul_34_17_n_9291 = ((mul_34_17_n_8653 & mul_34_17_n_8803) | ((mul_34_17_n_8653 & mul_34_17_n_8651)
    | (mul_34_17_n_8651 & mul_34_17_n_8803)));
 assign mul_34_17_n_9289 = ((mul_34_17_n_8754 & mul_34_17_n_8860) | ((mul_34_17_n_8754 & mul_34_17_n_8726)
    | (mul_34_17_n_8726 & mul_34_17_n_8860)));
 assign mul_34_17_n_9288 = ((mul_34_17_n_8756 & mul_34_17_n_8671) | ((mul_34_17_n_8756 & mul_34_17_n_8757)
    | (mul_34_17_n_8757 & mul_34_17_n_8671)));
 assign mul_34_17_n_9287 = ((mul_34_17_n_8770 & mul_34_17_n_269) | ((mul_34_17_n_8770 & mul_34_17_n_8546)
    | (mul_34_17_n_8546 & mul_34_17_n_269)));
 assign mul_34_17_n_9286 = ((mul_34_17_n_8794 & mul_34_17_n_8864) | ((mul_34_17_n_8794 & mul_34_17_n_8795)
    | (mul_34_17_n_8795 & mul_34_17_n_8864)));
 assign mul_34_17_n_9285 = ((mul_34_17_n_7941 & mul_34_17_n_8881) | ((mul_34_17_n_7941 & mul_34_17_n_7798)
    | (mul_34_17_n_7798 & mul_34_17_n_8881)));
 assign mul_34_17_n_9231 = ~(mul_34_17_n_236 | mul_34_17_n_8791);
 assign mul_34_17_n_9230 = ~(mul_34_17_n_9036 | mul_34_17_n_8790);
 assign mul_34_17_n_9284 = ((mul_34_17_n_8607 & mul_34_17_n_8566) | ((mul_34_17_n_8607 & mul_34_17_n_8332)
    | (mul_34_17_n_8332 & mul_34_17_n_8566)));
 assign mul_34_17_n_9283 = ((mul_34_17_n_8624 & mul_34_17_n_8491) | ((mul_34_17_n_8624 & mul_34_17_n_8498)
    | (mul_34_17_n_8498 & mul_34_17_n_8491)));
 assign mul_34_17_n_9281 = ((mul_34_17_n_8797 & mul_34_17_n_8935) | ((mul_34_17_n_8797 & mul_34_17_n_8796)
    | (mul_34_17_n_8796 & mul_34_17_n_8935)));
 assign mul_34_17_n_9280 = ((mul_34_17_n_8755 & mul_34_17_n_8943) | ((mul_34_17_n_8755 & mul_34_17_n_8532)
    | (mul_34_17_n_8532 & mul_34_17_n_8943)));
 assign mul_34_17_n_9279 = ~(mul_34_17_n_8882 ^ mul_34_17_n_8557);
 assign mul_34_17_n_9278 = ((mul_34_17_n_8389 & mul_34_17_n_8868) | ((mul_34_17_n_8389 & mul_34_17_n_8254)
    | (mul_34_17_n_8254 & mul_34_17_n_8868)));
 assign mul_34_17_n_9277 = ((mul_34_17_n_8766 & mul_34_17_n_8782) | ((mul_34_17_n_8766 & mul_34_17_n_8252)
    | (mul_34_17_n_8252 & mul_34_17_n_8782)));
 assign mul_34_17_n_9276 = (mul_34_17_n_11619 ^ mul_34_17_n_8745);
 assign mul_34_17_n_9275 = ((mul_34_17_n_8749 & mul_34_17_n_8563) | ((mul_34_17_n_8749 & mul_34_17_n_8359)
    | (mul_34_17_n_8359 & mul_34_17_n_8563)));
 assign mul_34_17_n_9274 = ((mul_34_17_n_8600 & mul_34_17_n_8948) | ((mul_34_17_n_8600 & mul_34_17_n_8719)
    | (mul_34_17_n_8719 & mul_34_17_n_8948)));
 assign mul_34_17_n_9273 = ~(mul_34_17_n_8860 ^ mul_34_17_n_251);
 assign mul_34_17_n_9272 = ((mul_34_17_n_8617 & mul_34_17_n_8674) | ((mul_34_17_n_8617 & mul_34_17_n_8232)
    | (mul_34_17_n_8232 & mul_34_17_n_8674)));
 assign mul_34_17_n_9271 = ((mul_34_17_n_8598 & mul_34_17_n_8407) | ((mul_34_17_n_8598 & mul_34_17_n_8008)
    | (mul_34_17_n_8008 & mul_34_17_n_8407)));
 assign mul_34_17_n_9270 = ~(mul_34_17_n_8885 ^ mul_34_17_n_8419);
 assign mul_34_17_n_9269 = ~((mul_34_17_n_8701 & mul_34_17_n_8562) | (mul_34_17_n_8905 & mul_34_17_n_8220));
 assign mul_34_17_n_9268 = ~(mul_34_17_n_8921 ^ mul_34_17_n_8325);
 assign mul_34_17_n_9267 = ((mul_34_17_n_8769 & mul_34_17_n_8863) | ((mul_34_17_n_8769 & mul_34_17_n_8510)
    | (mul_34_17_n_8510 & mul_34_17_n_8863)));
 assign mul_34_17_n_9266 = ~(mul_34_17_n_8573 ^ (mul_34_17_n_8269 ^ (mul_34_17_n_8572 ^ mul_34_17_n_7915)));
 assign mul_34_17_n_9265 = ((mul_34_17_n_8744 & mul_34_17_n_8938) | ((mul_34_17_n_8744 & mul_34_17_n_8537)
    | (mul_34_17_n_8537 & mul_34_17_n_8938)));
 assign mul_34_17_n_9263 = ((mul_34_17_n_8664 & mul_34_17_n_8682) | ((mul_34_17_n_8664 & mul_34_17_n_8346)
    | (mul_34_17_n_8346 & mul_34_17_n_8682)));
 assign mul_34_17_n_9262 = ((mul_34_17_n_8746 & mul_34_17_n_8734) | ((mul_34_17_n_8746 & mul_34_17_n_8605)
    | (mul_34_17_n_8605 & mul_34_17_n_8734)));
 assign mul_34_17_n_9261 = ((mul_34_17_n_8623 & mul_34_17_n_235) | (mul_34_17_n_8902 & mul_34_17_n_8677));
 assign mul_34_17_n_9260 = ((mul_34_17_n_11366 & mul_34_17_n_8789) | ((mul_34_17_n_11366 & mul_34_17_n_8743)
    | (mul_34_17_n_8743 & mul_34_17_n_8789)));
 assign mul_34_17_n_9225 = ~mul_34_17_n_9224;
 assign mul_34_17_n_9212 = ~mul_34_17_n_9211;
 assign mul_34_17_n_9198 = ~mul_34_17_n_9197;
 assign mul_34_17_n_9181 = ~mul_34_17_n_9182;
 assign mul_34_17_n_9175 = ~mul_34_17_n_9174;
 assign mul_34_17_n_9169 = ~mul_34_17_n_11326;
 assign mul_34_17_n_9154 = ~(mul_34_17_n_8835 ^ mul_34_17_n_8595);
 assign mul_34_17_n_9153 = (mul_34_17_n_8855 ^ mul_34_17_n_8495);
 assign mul_34_17_n_9229 = (mul_34_17_n_8619 ^ mul_34_17_n_8845);
 assign mul_34_17_n_9152 = (mul_34_17_n_11621 ^ mul_34_17_n_8841);
 assign mul_34_17_n_9228 = ~(mul_34_17_n_8823 ^ mul_34_17_n_8240);
 assign mul_34_17_n_9227 = ((mul_34_17_n_8591 & mul_34_17_n_8842) | ((mul_34_17_n_8591 & mul_34_17_n_8603)
    | (mul_34_17_n_8603 & mul_34_17_n_8842)));
 assign mul_34_17_n_9226 = ~(mul_34_17_n_8405 ^ (mul_34_17_n_8249 ^ (mul_34_17_n_8162 ^ mul_34_17_n_7781)));
 assign mul_34_17_n_9224 = ((mul_34_17_n_8649 & mul_34_17_n_8406) | ((mul_34_17_n_8649 & mul_34_17_n_8530)
    | (mul_34_17_n_8530 & mul_34_17_n_8406)));
 assign mul_34_17_n_9151 = (mul_34_17_n_8853 ^ mul_34_17_n_8650);
 assign mul_34_17_n_9150 = (mul_34_17_n_244 ^ mul_34_17_n_8625);
 assign mul_34_17_n_9223 = ((mul_34_17_n_8652 & mul_34_17_n_8666) | ((mul_34_17_n_8652 & mul_34_17_n_8538)
    | (mul_34_17_n_8538 & mul_34_17_n_8666)));
 assign mul_34_17_n_9222 = ((mul_34_17_n_8518 & mul_34_17_n_8941) | ((mul_34_17_n_8518 & mul_34_17_n_8540)
    | (mul_34_17_n_8540 & mul_34_17_n_8941)));
 assign mul_34_17_n_9221 = (mul_34_17_n_8863 ^ mul_34_17_n_8510);
 assign mul_34_17_n_9220 = ~(mul_34_17_n_8808 ^ mul_34_17_n_8494);
 assign mul_34_17_n_9149 = ~(mul_34_17_n_8424 ^ (mul_34_17_n_7890 ^ (mul_34_17_n_8169 ^ mul_34_17_n_7515)));
 assign mul_34_17_n_9148 = ~(mul_34_17_n_8873 ^ mul_34_17_n_8248);
 assign mul_34_17_n_9147 = ~(mul_34_17_n_8598 ^ mul_34_17_n_8850);
 assign mul_34_17_n_9219 = ~(mul_34_17_n_8886 ^ mul_34_17_n_8402);
 assign mul_34_17_n_9218 = (mul_34_17_n_259 ^ mul_34_17_n_256);
 assign mul_34_17_n_9146 = (mul_34_17_n_8874 ^ mul_34_17_n_8633);
 assign mul_34_17_n_9217 = (mul_34_17_n_8923 ^ mul_34_17_n_8640);
 assign mul_34_17_n_9145 = ~(mul_34_17_n_8868 ^ mul_34_17_n_8389);
 assign mul_34_17_n_9144 = (mul_34_17_n_8876 ^ mul_34_17_n_8381);
 assign mul_34_17_n_9143 = (mul_34_17_n_8632 ^ mul_34_17_n_11336);
 assign mul_34_17_n_9216 = ((mul_34_17_n_8731 & mul_34_17_n_8918) | ((mul_34_17_n_8731 & mul_34_17_n_8553)
    | (mul_34_17_n_8553 & mul_34_17_n_8918)));
 assign mul_34_17_n_9142 = (mul_34_17_n_8866 ^ mul_34_17_n_8933);
 assign mul_34_17_n_9141 = (mul_34_17_n_8949 ^ mul_34_17_n_8930);
 assign mul_34_17_n_9140 = ~((mul_34_17_n_7326 & (~mul_34_17_n_7341 & ~mul_34_17_n_8889)) | ((mul_34_17_n_7325
    & (mul_34_17_n_7341 & ~mul_34_17_n_8889)) | (mul_34_17_n_7960 & mul_34_17_n_8889)));
 assign mul_34_17_n_9215 = ~(mul_34_17_n_8897 ^ mul_34_17_n_11623);
 assign mul_34_17_n_9214 = ((mul_34_17_n_8648 & mul_34_17_n_8686) | ((mul_34_17_n_8648 & mul_34_17_n_8379)
    | (mul_34_17_n_8379 & mul_34_17_n_8686)));
 assign mul_34_17_n_9213 = ((mul_34_17_n_8641 & mul_34_17_n_8875) | ((mul_34_17_n_8641 & mul_34_17_n_8339)
    | (mul_34_17_n_8339 & mul_34_17_n_8875)));
 assign mul_34_17_n_9211 = ((mul_34_17_n_8615 & mul_34_17_n_8404) | ((mul_34_17_n_8615 & mul_34_17_n_8250)
    | (mul_34_17_n_8250 & mul_34_17_n_8404)));
 assign mul_34_17_n_9210 = ((mul_34_17_n_364 & mul_34_17_n_8556) | (mul_34_17_n_8904 & mul_34_17_n_8206));
 assign mul_34_17_n_9209 = ~(mul_34_17_n_8383 ^ (mul_34_17_n_8266 ^ (mul_34_17_n_7940 ^ mul_34_17_n_7103)));
 assign mul_34_17_n_9208 = ~(mul_34_17_n_8891 ^ mul_34_17_n_8497);
 assign mul_34_17_n_9207 = ~(mul_34_17_n_8844 ^ mul_34_17_n_8128);
 assign mul_34_17_n_9206 = ((mul_34_17_n_11354 & mul_34_17_n_8680) | ((mul_34_17_n_11354 & mul_34_17_n_255)
    | (mul_34_17_n_255 & mul_34_17_n_8680)));
 assign mul_34_17_n_9205 = ((mul_34_17_n_8670 & mul_34_17_n_8611) | ((mul_34_17_n_8670 & mul_34_17_n_8593)
    | (mul_34_17_n_8593 & mul_34_17_n_8611)));
 assign mul_34_17_n_9204 = ((mul_34_17_n_8662 & mul_34_17_n_8835) | ((mul_34_17_n_8662 & mul_34_17_n_8594)
    | (mul_34_17_n_8594 & mul_34_17_n_8835)));
 assign mul_34_17_n_9203 = ~((mul_34_17_n_7427 & (~mul_34_17_n_8367 & ~mul_34_17_n_8445)) | ((mul_34_17_n_7428
    & (mul_34_17_n_8367 & ~mul_34_17_n_8445)) | (mul_34_17_n_8881 & mul_34_17_n_8445)));
 assign mul_34_17_n_9202 = ((mul_34_17_n_8747 & mul_34_17_n_8786) | ((mul_34_17_n_8747 & mul_34_17_n_8748)
    | (mul_34_17_n_8748 & mul_34_17_n_8786)));
 assign mul_34_17_n_9200 = ~(mul_34_17_n_8895 ^ mul_34_17_n_8504);
 assign mul_34_17_n_9199 = ~(mul_34_17_n_8819 ^ mul_34_17_n_11360);
 assign mul_34_17_n_9197 = ~(mul_34_17_n_8818 ^ mul_34_17_n_8776);
 assign mul_34_17_n_9196 = ((mul_34_17_n_8759 & mul_34_17_n_8945) | ((mul_34_17_n_8759 & mul_34_17_n_8758)
    | (mul_34_17_n_8758 & mul_34_17_n_8945)));
 assign mul_34_17_n_9195 = ~(mul_34_17_n_8807 ^ mul_34_17_n_8366);
 assign mul_34_17_n_9194 = (mul_34_17_n_8843 ^ mul_34_17_n_8867);
 assign mul_34_17_n_9193 = ~(mul_34_17_n_8809 ^ mul_34_17_n_8242);
 assign mul_34_17_n_9192 = ((mul_34_17_n_8771 & mul_34_17_n_8561) | ((mul_34_17_n_8771 & mul_34_17_n_8500)
    | (mul_34_17_n_8500 & mul_34_17_n_8561)));
 assign mul_34_17_n_9191 = ~(mul_34_17_n_8806 ^ mul_34_17_n_8344);
 assign mul_34_17_n_9190 = ((mul_34_17_n_8638 & mul_34_17_n_8417) | ((mul_34_17_n_8638 & mul_34_17_n_8639)
    | (mul_34_17_n_8639 & mul_34_17_n_8417)));
 assign mul_34_17_n_9189 = ~(mul_34_17_n_8813 ^ mul_34_17_n_8336);
 assign mul_34_17_n_9188 = ((mul_34_17_n_8362 & mul_34_17_n_8937) | ((mul_34_17_n_8362 & mul_34_17_n_8356)
    | (mul_34_17_n_8356 & mul_34_17_n_8937)));
 assign mul_34_17_n_9187 = ~(mul_34_17_n_8820 ^ mul_34_17_n_8410);
 assign mul_34_17_n_9186 = ~(mul_34_17_n_8810 ^ mul_34_17_n_8528);
 assign mul_34_17_n_9185 = (mul_34_17_n_11344 ^ mul_34_17_n_8631);
 assign mul_34_17_n_9184 = ~(mul_34_17_n_8812 ^ mul_34_17_n_11372);
 assign mul_34_17_n_9183 = ((mul_34_17_n_8576 & mul_34_17_n_8578) | ((mul_34_17_n_8576 & mul_34_17_n_8370)
    | (mul_34_17_n_8370 & mul_34_17_n_8578)));
 assign mul_34_17_n_9182 = (mul_34_17_n_8880 ^ mul_34_17_n_8385);
 assign mul_34_17_n_9180 = ((mul_34_17_n_8661 & mul_34_17_n_11356) | ((mul_34_17_n_8661 & mul_34_17_n_8657)
    | (mul_34_17_n_8657 & mul_34_17_n_11356)));
 assign mul_34_17_n_9179 = ~((mul_34_17_n_7979 & (~mul_34_17_n_8489 & ~mul_34_17_n_8610)) | ((mul_34_17_n_7980
    & (mul_34_17_n_8489 & ~mul_34_17_n_8610)) | (mul_34_17_n_8901 & mul_34_17_n_8610)));
 assign mul_34_17_n_9178 = ~(mul_34_17_n_8814 ^ mul_34_17_n_8365);
 assign mul_34_17_n_9177 = ((mul_34_17_n_246 & mul_34_17_n_8916) | ((mul_34_17_n_246 & mul_34_17_n_8533)
    | (mul_34_17_n_8533 & mul_34_17_n_8916)));
 assign mul_34_17_n_9176 = ~(mul_34_17_n_8815 ^ mul_34_17_n_8503);
 assign mul_34_17_n_9174 = ((mul_34_17_n_8612 & mul_34_17_n_8870) | ((mul_34_17_n_8612 & mul_34_17_n_8333)
    | (mul_34_17_n_8333 & mul_34_17_n_8870)));
 assign mul_34_17_n_9173 = ((mul_34_17_n_8620 & mul_34_17_n_8330) | ((mul_34_17_n_8620 & mul_34_17_n_8328)
    | (mul_34_17_n_8328 & mul_34_17_n_8330)));
 assign mul_34_17_n_9172 = ~(mul_34_17_n_8821 ^ mul_34_17_n_8376);
 assign mul_34_17_n_9171 = ((mul_34_17_n_8658 & mul_34_17_n_8939) | ((mul_34_17_n_8658 & mul_34_17_n_8138)
    | (mul_34_17_n_8138 & mul_34_17_n_8939)));
 assign mul_34_17_n_9170 = (mul_34_17_n_230 ^ mul_34_17_n_8382);
 assign mul_34_17_n_9167 = ~((mul_34_17_n_8329 & (~mul_34_17_n_8330 & ~mul_34_17_n_8620)) | ((mul_34_17_n_8328
    & (mul_34_17_n_8330 & ~mul_34_17_n_8620)) | (mul_34_17_n_8825 & mul_34_17_n_8620)));
 assign mul_34_17_n_9166 = ((mul_34_17_n_8613 & mul_34_17_n_11352) | ((mul_34_17_n_8613 & mul_34_17_n_8663)
    | (mul_34_17_n_8663 & mul_34_17_n_11352)));
 assign mul_34_17_n_9164 = ((mul_34_17_n_8587 & mul_34_17_n_7928) | (mul_34_17_n_8908 & mul_34_17_n_7637));
 assign mul_34_17_n_9163 = ((mul_34_17_n_8654 & mul_34_17_n_11374) | ((mul_34_17_n_8654 & mul_34_17_n_8375)
    | (mul_34_17_n_8375 & mul_34_17_n_11374)));
 assign mul_34_17_n_9162 = ~(mul_34_17_n_8816 ^ mul_34_17_n_8386);
 assign mul_34_17_n_9160 = ((mul_34_17_n_8630 & mul_34_17_n_8877) | ((mul_34_17_n_8630 & mul_34_17_n_8629)
    | (mul_34_17_n_8629 & mul_34_17_n_8877)));
 assign mul_34_17_n_9159 = (mul_34_17_n_8952 ^ mul_34_17_n_8409);
 assign mul_34_17_n_9158 = ((mul_34_17_n_8577 & mul_34_17_n_8684) | ((mul_34_17_n_8577 & mul_34_17_n_8282)
    | (mul_34_17_n_8282 & mul_34_17_n_8684)));
 assign mul_34_17_n_9139 = ~mul_34_17_n_9074;
 assign mul_34_17_n_9133 = ~mul_34_17_n_9132;
 assign mul_34_17_n_9131 = ~mul_34_17_n_9047;
 assign mul_34_17_n_9127 = ~mul_34_17_n_9126;
 assign mul_34_17_n_9122 = ~mul_34_17_n_9121;
 assign mul_34_17_n_9116 = ~mul_34_17_n_9117;
 assign mul_34_17_n_9106 = ~mul_34_17_n_9107;
 assign mul_34_17_n_9096 = ~mul_34_17_n_9095;
 assign mul_34_17_n_9091 = ~mul_34_17_n_9092;
 assign mul_34_17_n_9087 = ~(mul_34_17_n_8906 | mul_34_17_n_8405);
 assign mul_34_17_n_9086 = (mul_34_17_n_8770 ^ mul_34_17_n_8546);
 assign mul_34_17_n_9084 = ~(mul_34_17_n_8844 & mul_34_17_n_8128);
 assign mul_34_17_n_9083 = ~(mul_34_17_n_8844 | mul_34_17_n_8128);
 assign mul_34_17_n_9082 = ~(mul_34_17_n_8921 & mul_34_17_n_8325);
 assign mul_34_17_n_9081 = ~(mul_34_17_n_8921 | mul_34_17_n_8325);
 assign mul_34_17_n_9080 = ~(mul_34_17_n_8653 ^ mul_34_17_n_8651);
 assign mul_34_17_n_9079 = ~(mul_34_17_n_8688 ^ mul_34_17_n_8428);
 assign mul_34_17_n_9078 = ~(mul_34_17_n_8848 & mul_34_17_n_8324);
 assign mul_34_17_n_9077 = ~(mul_34_17_n_259 & mul_34_17_n_8660);
 assign mul_34_17_n_9076 = ~(mul_34_17_n_8856 & mul_34_17_n_256);
 assign mul_34_17_n_9075 = ~(mul_34_17_n_8848 | mul_34_17_n_8324);
 assign mul_34_17_n_9074 = ~(mul_34_17_n_259 | mul_34_17_n_256);
 assign mul_34_17_n_9073 = ((mul_34_17_n_7902 & mul_34_17_n_7751) | (mul_34_17_n_8799 & mul_34_17_n_8280));
 assign mul_34_17_n_9072 = ~(mul_34_17_n_8689 ^ mul_34_17_n_8274);
 assign mul_34_17_n_9071 = ~(mul_34_17_n_8946 & mul_34_17_n_8431);
 assign mul_34_17_n_9069 = ~(mul_34_17_n_259 & mul_34_17_n_256);
 assign mul_34_17_n_9068 = ~(mul_34_17_n_8720 ^ mul_34_17_n_8599);
 assign mul_34_17_n_9067 = ~(mul_34_17_n_8276 ^ (mul_34_17_n_7788 ^ (mul_34_17_n_8069 ^ mul_34_17_n_7696)));
 assign mul_34_17_n_9066 = ~(mul_34_17_n_8060 ^ (mul_34_17_n_8166 ^ (mul_34_17_n_7936 ^ mul_34_17_n_7350)));
 assign mul_34_17_n_9065 = ~(mul_34_17_n_8855 & mul_34_17_n_8495);
 assign mul_34_17_n_9064 = ~(mul_34_17_n_8687 ^ mul_34_17_n_8425);
 assign mul_34_17_n_9063 = ~(mul_34_17_n_8797 ^ mul_34_17_n_8796);
 assign mul_34_17_n_9062 = ~(mul_34_17_n_8896 & mul_34_17_n_8272);
 assign mul_34_17_n_9061 = ~(mul_34_17_n_8802 ^ mul_34_17_n_11350);
 assign mul_34_17_n_9060 = (mul_34_17_n_8751 ^ mul_34_17_n_8753);
 assign mul_34_17_n_9059 = (mul_34_17_n_8747 ^ mul_34_17_n_8748);
 assign mul_34_17_n_9058 = (mul_34_17_n_8757 ^ mul_34_17_n_8671);
 assign mul_34_17_n_9057 = ~(mul_34_17_n_8783 ^ mul_34_17_n_8520);
 assign mul_34_17_n_9056 = (mul_34_17_n_8771 ^ mul_34_17_n_8561);
 assign mul_34_17_n_9138 = ~(mul_34_17_n_8659 ^ mul_34_17_n_8373);
 assign mul_34_17_n_9137 = ~(mul_34_17_n_8947 | mul_34_17_n_8430);
 assign mul_34_17_n_9055 = (mul_34_17_n_8763 ^ mul_34_17_n_8762);
 assign mul_34_17_n_9054 = ~(mul_34_17_n_8668 ^ mul_34_17_n_8501);
 assign mul_34_17_n_9053 = ~(mul_34_17_n_8794 ^ mul_34_17_n_8795);
 assign mul_34_17_n_9052 = ~(mul_34_17_n_11358 ^ mul_34_17_n_8394);
 assign mul_34_17_n_9051 = ~(mul_34_17_n_8623 ^ mul_34_17_n_8673);
 assign mul_34_17_n_9136 = ~(mul_34_17_n_8855 | mul_34_17_n_8495);
 assign mul_34_17_n_9050 = (mul_34_17_n_8755 ^ mul_34_17_n_8532);
 assign mul_34_17_n_9049 = ~(mul_34_17_n_8787 ^ mul_34_17_n_8515);
 assign mul_34_17_n_9048 = (mul_34_17_n_8563 ^ mul_34_17_n_8749);
 assign mul_34_17_n_9134 = ((mul_34_17_n_8338 & mul_34_17_n_8402) | ((mul_34_17_n_8338 & mul_34_17_n_8509)
    | (mul_34_17_n_8509 & mul_34_17_n_8402)));
 assign mul_34_17_n_9132 = ~(mul_34_17_n_11334 | mul_34_17_n_8804);
 assign mul_34_17_n_9047 = ~(mul_34_17_n_8879 & mul_34_17_n_8423);
 assign mul_34_17_n_9130 = ((mul_34_17_n_11378 & mul_34_17_n_8777) | ((mul_34_17_n_11378 & mul_34_17_n_8525)
    | (mul_34_17_n_8525 & mul_34_17_n_8777)));
 assign mul_34_17_n_9129 = ((mul_34_17_n_8511 & mul_34_17_n_8262) | ((mul_34_17_n_8511 & mul_34_17_n_11400)
    | (mul_34_17_n_11400 & mul_34_17_n_8262)));
 assign mul_34_17_n_9128 = ~((mul_34_17_n_371 & mul_34_17_n_8049) | (mul_34_17_n_8715 & mul_34_17_n_7659));
 assign mul_34_17_n_9126 = ~(mul_34_17_n_8691 ^ mul_34_17_n_8234);
 assign mul_34_17_n_9125 = ((mul_34_17_n_8451 & mul_34_17_n_8064) | (mul_34_17_n_8700 & mul_34_17_n_7663));
 assign mul_34_17_n_9124 = ((mul_34_17_n_8454 & mul_34_17_n_8559) | (mul_34_17_n_8714 & mul_34_17_n_8216));
 assign mul_34_17_n_9123 = ((mul_34_17_n_8354 & mul_34_17_n_8420) | ((mul_34_17_n_8354 & mul_34_17_n_8242)
    | (mul_34_17_n_8242 & mul_34_17_n_8420)));
 assign mul_34_17_n_9121 = ((mul_34_17_n_8388 & mul_34_17_n_11360) | ((mul_34_17_n_8388 & mul_34_17_n_8527)
    | (mul_34_17_n_8527 & mul_34_17_n_11360)));
 assign mul_34_17_n_9120 = ((mul_34_17_n_8341 & mul_34_17_n_8558) | ((mul_34_17_n_8341 & mul_34_17_n_8013)
    | (mul_34_17_n_8013 & mul_34_17_n_8558)));
 assign mul_34_17_n_9119 = ((mul_34_17_n_8374 & mul_34_17_n_7926) | ((mul_34_17_n_8374 & mul_34_17_n_11456)
    | (mul_34_17_n_11456 & mul_34_17_n_7926)));
 assign mul_34_17_n_9118 = ((mul_34_17_n_8485 & mul_34_17_n_8227) | ((mul_34_17_n_8485 & mul_34_17_n_8524)
    | (mul_34_17_n_8524 & mul_34_17_n_8227)));
 assign mul_34_17_n_9117 = ((mul_34_17_n_8502 & mul_34_17_n_8669) | ((mul_34_17_n_8502 & mul_34_17_n_8512)
    | (mul_34_17_n_8512 & mul_34_17_n_8669)));
 assign mul_34_17_n_9115 = ((mul_34_17_n_8545 & mul_34_17_n_8780) | ((mul_34_17_n_8545 & mul_34_17_n_8032)
    | (mul_34_17_n_8032 & mul_34_17_n_8780)));
 assign mul_34_17_n_9114 = ((mul_34_17_n_8516 & mul_34_17_n_8157) | ((mul_34_17_n_8516 & mul_34_17_n_232)
    | (mul_34_17_n_232 & mul_34_17_n_8157)));
 assign mul_34_17_n_9113 = ~(mul_34_17_n_8784 ^ mul_34_17_n_8535);
 assign mul_34_17_n_9112 = ((mul_34_17_n_8497 & mul_34_17_n_11376) | ((mul_34_17_n_8497 & mul_34_17_n_11454)
    | (mul_34_17_n_11454 & mul_34_17_n_11376)));
 assign mul_34_17_n_9111 = ((mul_34_17_n_8486 & mul_34_17_n_8256) | ((mul_34_17_n_8486 & mul_34_17_n_7898)
    | (mul_34_17_n_7898 & mul_34_17_n_8256)));
 assign mul_34_17_n_9110 = ((mul_34_17_n_8342 & mul_34_17_n_8259) | ((mul_34_17_n_8342 & mul_34_17_n_8344)
    | (mul_34_17_n_8344 & mul_34_17_n_8259)));
 assign mul_34_17_n_9109 = ((mul_34_17_n_8531 & mul_34_17_n_8403) | ((mul_34_17_n_8531 & mul_34_17_n_8536)
    | (mul_34_17_n_8536 & mul_34_17_n_8403)));
 assign mul_34_17_n_9108 = ((mul_34_17_n_8363 & mul_34_17_n_8672) | ((mul_34_17_n_8363 & mul_34_17_n_8505)
    | (mul_34_17_n_8505 & mul_34_17_n_8672)));
 assign mul_34_17_n_9107 = ((mul_34_17_n_11380 & mul_34_17_n_11384) | ((mul_34_17_n_11380 & mul_34_17_n_8504)
    | (mul_34_17_n_8504 & mul_34_17_n_11384)));
 assign mul_34_17_n_9105 = ((mul_34_17_n_8547 & mul_34_17_n_8062) | ((mul_34_17_n_8547 & mul_34_17_n_8245)
    | (mul_34_17_n_8245 & mul_34_17_n_8062)));
 assign mul_34_17_n_9104 = ((mul_34_17_n_8327 & mul_34_17_n_8152) | ((mul_34_17_n_8327 & mul_34_17_n_8236)
    | (mul_34_17_n_8236 & mul_34_17_n_8152)));
 assign mul_34_17_n_9102 = ((mul_34_17_n_8515 & mul_34_17_n_8788) | ((mul_34_17_n_8515 & mul_34_17_n_8550)
    | (mul_34_17_n_8550 & mul_34_17_n_8788)));
 assign mul_34_17_n_9101 = ~(mul_34_17_n_8696 ^ mul_34_17_n_8547);
 assign mul_34_17_n_9100 = ((mul_34_17_n_8556 & mul_34_17_n_8223) | ((mul_34_17_n_8556 & mul_34_17_n_7668)
    | (mul_34_17_n_7668 & mul_34_17_n_8223)));
 assign mul_34_17_n_9099 = ((mul_34_17_n_8340 & mul_34_17_n_11382) | ((mul_34_17_n_8340 & mul_34_17_n_8023)
    | (mul_34_17_n_8023 & mul_34_17_n_11382)));
 assign mul_34_17_n_9098 = ((mul_34_17_n_8707 & mul_34_17_n_8469) | (mul_34_17_n_8711 & mul_34_17_n_234));
 assign mul_34_17_n_9097 = (mul_34_17_n_8568 ^ mul_34_17_n_8750);
 assign mul_34_17_n_9095 = ((mul_34_17_n_234 & mul_34_17_n_8231) | ((mul_34_17_n_234 & mul_34_17_n_228)
    | (mul_34_17_n_228 & mul_34_17_n_8231)));
 assign mul_34_17_n_9094 = ~(mul_34_17_n_8695 ^ mul_34_17_n_8555);
 assign mul_34_17_n_9093 = ((mul_34_17_n_8503 & mul_34_17_n_8554) | ((mul_34_17_n_8503 & mul_34_17_n_8506)
    | (mul_34_17_n_8506 & mul_34_17_n_8554)));
 assign mul_34_17_n_9092 = ((mul_34_17_n_231 & mul_34_17_n_8557) | ((mul_34_17_n_231 & mul_34_17_n_8534)
    | (mul_34_17_n_8534 & mul_34_17_n_8557)));
 assign mul_34_17_n_9090 = ((mul_34_17_n_8528 & mul_34_17_n_8418) | ((mul_34_17_n_8528 & mul_34_17_n_7899)
    | (mul_34_17_n_7899 & mul_34_17_n_8418)));
 assign mul_34_17_n_9089 = ~((mul_34_17_n_8459 & mul_34_17_n_8054) | (mul_34_17_n_8713 & mul_34_17_n_7654));
 assign mul_34_17_n_9088 = ((mul_34_17_n_8521 & mul_34_17_n_8783) | ((mul_34_17_n_8521 & mul_34_17_n_8529)
    | (mul_34_17_n_8529 & mul_34_17_n_8783)));
 assign mul_34_17_n_9036 = ~mul_34_17_n_236;
 assign mul_34_17_n_9034 = ~mul_34_17_n_275;
 assign mul_34_17_n_9010 = ~mul_34_17_n_9009;
 assign mul_34_17_n_9001 = ~mul_34_17_n_9000;
 assign mul_34_17_n_8997 = ~mul_34_17_n_8996;
 assign mul_34_17_n_8989 = ~mul_34_17_n_8988;
 assign mul_34_17_n_8981 = ~(mul_34_17_n_8734 ^ mul_34_17_n_11368);
 assign mul_34_17_n_8976 = ~(mul_34_17_n_8172 ^ (mul_34_17_n_202 ^ (mul_34_17_n_8173 ^ mul_34_17_n_7085)));
 assign mul_34_17_n_8975 = ~(mul_34_17_n_8167 ^ (mul_34_17_n_11637 ^ (mul_34_17_n_8159 ^ mul_34_17_n_7592)));
 assign mul_34_17_n_8974 = ~((mul_34_17_n_8314 | mul_34_17_n_7980) & (mul_34_17_n_8610 | mul_34_17_n_8693));
 assign mul_34_17_n_9046 = ~(mul_34_17_n_8642 ^ mul_34_17_n_8327);
 assign mul_34_17_n_9045 = ((mul_34_17_n_8348 & mul_34_17_n_8268) | ((mul_34_17_n_8348 & mul_34_17_n_8513)
    | (mul_34_17_n_8513 & mul_34_17_n_8268)));
 assign mul_34_17_n_9044 = ((mul_34_17_n_8542 & mul_34_17_n_8551) | ((mul_34_17_n_8542 & mul_34_17_n_8523)
    | (mul_34_17_n_8523 & mul_34_17_n_8551)));
 assign mul_34_17_n_8971 = (mul_34_17_n_8648 ^ mul_34_17_n_8686);
 assign mul_34_17_n_8970 = (mul_34_17_n_8617 ^ mul_34_17_n_8674);
 assign mul_34_17_n_9043 = (mul_34_17_n_11354 ^ mul_34_17_n_255);
 assign mul_34_17_n_8969 = (mul_34_17_n_8417 ^ mul_34_17_n_8639);
 assign mul_34_17_n_8968 = (mul_34_17_n_11352 ^ mul_34_17_n_8613);
 assign mul_34_17_n_8967 = ~(mul_34_17_n_8607 ^ mul_34_17_n_8331);
 assign mul_34_17_n_9042 = (mul_34_17_n_11374 ^ mul_34_17_n_8654);
 assign mul_34_17_n_8966 = (mul_34_17_n_8538 ^ mul_34_17_n_8652);
 assign mul_34_17_n_9041 = ((mul_34_17_n_226 & mul_34_17_n_8129) | ((mul_34_17_n_226 & mul_34_17_n_7422)
    | (mul_34_17_n_7422 & mul_34_17_n_8129)));
 assign mul_34_17_n_8965 = (mul_34_17_n_8672 ^ mul_34_17_n_8505);
 assign mul_34_17_n_9040 = ((mul_34_17_n_8384 & mul_34_17_n_8415) | ((mul_34_17_n_8384 & mul_34_17_n_8385)
    | (mul_34_17_n_8385 & mul_34_17_n_8415)));
 assign mul_34_17_n_9039 = ~(mul_34_17_n_8580 ^ mul_34_17_n_8390);
 assign mul_34_17_n_8964 = (mul_34_17_n_8743 ^ mul_34_17_n_11366);
 assign mul_34_17_n_8963 = ~(mul_34_17_n_8641 ^ mul_34_17_n_8339);
 assign mul_34_17_n_8962 = (mul_34_17_n_8530 ^ mul_34_17_n_8649);
 assign mul_34_17_n_8961 = (mul_34_17_n_8630 ^ mul_34_17_n_8629);
 assign mul_34_17_n_8960 = (mul_34_17_n_8621 ^ mul_34_17_n_8247);
 assign mul_34_17_n_9038 = ~(mul_34_17_n_8257 ^ mul_34_17_n_8694);
 assign mul_34_17_n_8959 = ~(mul_34_17_n_8675 ^ mul_34_17_n_8237);
 assign mul_34_17_n_8958 = ~(mul_34_17_n_8160 ^ (mul_34_17_n_8161 ^ (mul_34_17_n_7939 ^ mul_34_17_n_7383)));
 assign mul_34_17_n_8957 = (mul_34_17_n_8138 ^ mul_34_17_n_8658);
 assign mul_34_17_n_9037 = ((mul_34_17_n_8376 & mul_34_17_n_8158) | ((mul_34_17_n_8376 & mul_34_17_n_8377)
    | (mul_34_17_n_8377 & mul_34_17_n_8158)));
 assign mul_34_17_n_8956 = (mul_34_17_n_8150 ^ mul_34_17_n_8740);
 assign mul_34_17_n_8955 = ~(mul_34_17_n_8170 ^ (mul_34_17_n_7518 ^ (mul_34_17_n_8168 ^ mul_34_17_n_7567)));
 assign mul_34_17_n_8954 = (mul_34_17_n_8661 ^ mul_34_17_n_11356);
 assign mul_34_17_n_9035 = ((mul_34_17_n_8395 & mul_34_17_n_11358) | ((mul_34_17_n_8395 & mul_34_17_n_8393)
    | (mul_34_17_n_8393 & mul_34_17_n_11358)));
 assign mul_34_17_n_9033 = ((mul_34_17_n_8312 & mul_34_17_n_7931) | (mul_34_17_n_8710 & mul_34_17_n_7636));
 assign mul_34_17_n_9031 = ~(mul_34_17_n_8582 ^ mul_34_17_n_7754);
 assign mul_34_17_n_9030 = ((mul_34_17_n_366 & mul_34_17_n_7934) | (mul_34_17_n_8705 & mul_34_17_n_7617));
 assign mul_34_17_n_9029 = ((mul_34_17_n_8336 & mul_34_17_n_11625) | ((mul_34_17_n_8336 & mul_34_17_n_8398)
    | (mul_34_17_n_8398 & mul_34_17_n_11625)));
 assign mul_34_17_n_9028 = ((mul_34_17_n_365 & mul_34_17_n_7933) | (mul_34_17_n_8704 & mul_34_17_n_7615));
 assign mul_34_17_n_9027 = ((mul_34_17_n_8323 & mul_34_17_n_8266) | ((mul_34_17_n_8323 & mul_34_17_n_8383)
    | (mul_34_17_n_8383 & mul_34_17_n_8266)));
 assign mul_34_17_n_9026 = ((mul_34_17_n_8541 & mul_34_17_n_8776) | ((mul_34_17_n_8541 & mul_34_17_n_7860)
    | (mul_34_17_n_7860 & mul_34_17_n_8776)));
 assign mul_34_17_n_9025 = ((mul_34_17_n_370 & mul_34_17_n_8055) | (mul_34_17_n_8712 & mul_34_17_n_7648));
 assign mul_34_17_n_9024 = ~(mul_34_17_n_8146 ^ (mul_34_17_n_7519 ^ (mul_34_17_n_7942 ^ mul_34_17_n_7787)));
 assign mul_34_17_n_9023 = ~((mul_34_17_n_7862 & (~mul_34_17_n_7430 & ~mul_34_17_n_8579)) | ((mul_34_17_n_7861
    & (mul_34_17_n_7430 & ~mul_34_17_n_8579)) | (mul_34_17_n_8414 & mul_34_17_n_8579)));
 assign mul_34_17_n_9021 = ~((mul_34_17_n_7422 & (~mul_34_17_n_8129 & ~mul_34_17_n_226)) | ((mul_34_17_n_7421
    & (mul_34_17_n_8129 & ~mul_34_17_n_226)) | (mul_34_17_n_8585 & mul_34_17_n_226)));
 assign mul_34_17_n_9019 = ((mul_34_17_n_8413 & mul_34_17_n_7906) | ((mul_34_17_n_8413 & mul_34_17_n_8241)
    | (mul_34_17_n_8241 & mul_34_17_n_7906)));
 assign mul_34_17_n_9018 = ((mul_34_17_n_8335 & mul_34_17_n_8149) | ((mul_34_17_n_8335 & mul_34_17_n_7712)
    | (mul_34_17_n_7712 & mul_34_17_n_8149)));
 assign mul_34_17_n_9017 = ((mul_34_17_n_8366 & mul_34_17_n_8263) | ((mul_34_17_n_8366 & mul_34_17_n_8364)
    | (mul_34_17_n_8364 & mul_34_17_n_8263)));
 assign mul_34_17_n_9014 = ((mul_34_17_n_8365 & mul_34_17_n_8408) | ((mul_34_17_n_8365 & mul_34_17_n_8360)
    | (mul_34_17_n_8360 & mul_34_17_n_8408)));
 assign mul_34_17_n_9013 = ~(mul_34_17_n_8584 ^ mul_34_17_n_8334);
 assign mul_34_17_n_9012 = (mul_34_17_n_246 ^ mul_34_17_n_8533);
 assign mul_34_17_n_9011 = ((mul_34_17_n_8372 & mul_34_17_n_8411) | ((mul_34_17_n_8372 & mul_34_17_n_8240)
    | (mul_34_17_n_8240 & mul_34_17_n_8411)));
 assign mul_34_17_n_9009 = ((mul_34_17_n_8369 & mul_34_17_n_8676) | ((mul_34_17_n_8369 & mul_34_17_n_8237)
    | (mul_34_17_n_8237 & mul_34_17_n_8676)));
 assign mul_34_17_n_9007 = ~(mul_34_17_n_8581 ^ mul_34_17_n_8516);
 assign mul_34_17_n_9006 = ~(mul_34_17_n_8624 ^ mul_34_17_n_8498);
 assign mul_34_17_n_9005 = ((mul_34_17_n_8368 & mul_34_17_n_11372) | ((mul_34_17_n_8368 & mul_34_17_n_8009)
    | (mul_34_17_n_8009 & mul_34_17_n_11372)));
 assign mul_34_17_n_9004 = ((mul_34_17_n_8357 & mul_34_17_n_8560) | ((mul_34_17_n_8357 & mul_34_17_n_8358)
    | (mul_34_17_n_8358 & mul_34_17_n_8560)));
 assign mul_34_17_n_9003 = ((mul_34_17_n_8371 & mul_34_17_n_8416) | ((mul_34_17_n_8371 & mul_34_17_n_8127)
    | (mul_34_17_n_8127 & mul_34_17_n_8416)));
 assign mul_34_17_n_9002 = ((mul_34_17_n_8559 & mul_34_17_n_7996) | ((mul_34_17_n_8559 & mul_34_17_n_7842)
    | (mul_34_17_n_7842 & mul_34_17_n_7996)));
 assign mul_34_17_n_9000 = ((mul_34_17_n_8337 & mul_34_17_n_11623) | ((mul_34_17_n_8337 & mul_34_17_n_8380)
    | (mul_34_17_n_8380 & mul_34_17_n_11623)));
 assign mul_34_17_n_8999 = ((mul_34_17_n_8496 & mul_34_17_n_8552) | ((mul_34_17_n_8496 & mul_34_17_n_8325)
    | (mul_34_17_n_8325 & mul_34_17_n_8552)));
 assign mul_34_17_n_8998 = ~(mul_34_17_n_8690 ^ mul_34_17_n_8511);
 assign mul_34_17_n_8996 = ((mul_34_17_n_8281 & mul_34_17_n_8147) | ((mul_34_17_n_8281 & mul_34_17_n_7520)
    | (mul_34_17_n_7520 & mul_34_17_n_8147)));
 assign mul_34_17_n_8995 = ((mul_34_17_n_8391 & mul_34_17_n_11388) | ((mul_34_17_n_8391 & mul_34_17_n_8145)
    | (mul_34_17_n_8145 & mul_34_17_n_11388)));
 assign mul_34_17_n_8993 = ~((mul_34_17_n_164 & (~mul_34_17_n_8228 & ~mul_34_17_n_7716)) | ((mul_34_17_n_7987
    & (mul_34_17_n_8228 & ~mul_34_17_n_7716)) | (mul_34_17_n_8590 & mul_34_17_n_7716)));
 assign mul_34_17_n_8992 = ~((mul_34_17_n_180 & (~mul_34_17_n_8130 & ~mul_34_17_n_7454)) | ((mul_34_17_n_7836
    & (mul_34_17_n_8130 & ~mul_34_17_n_7454)) | (mul_34_17_n_8589 & mul_34_17_n_7454)));
 assign mul_34_17_n_8991 = ((mul_34_17_n_8343 & mul_34_17_n_11370) | ((mul_34_17_n_8343 & mul_34_17_n_8387)
    | (mul_34_17_n_8387 & mul_34_17_n_11370)));
 assign mul_34_17_n_8990 = ((mul_34_17_n_8519 & mul_34_17_n_8410) | ((mul_34_17_n_8519 & mul_34_17_n_227)
    | (mul_34_17_n_227 & mul_34_17_n_8410)));
 assign mul_34_17_n_8988 = ((mul_34_17_n_8535 & mul_34_17_n_8785) | ((mul_34_17_n_8535 & mul_34_17_n_8487)
    | (mul_34_17_n_8487 & mul_34_17_n_8785)));
 assign mul_34_17_n_8987 = ((mul_34_17_n_8494 & mul_34_17_n_8564) | ((mul_34_17_n_8494 & mul_34_17_n_8392)
    | (mul_34_17_n_8392 & mul_34_17_n_8564)));
 assign mul_34_17_n_8986 = ((mul_34_17_n_8499 & mul_34_17_n_8775) | ((mul_34_17_n_8499 & mul_34_17_n_8355)
    | (mul_34_17_n_8355 & mul_34_17_n_8775)));
 assign mul_34_17_n_8985 = ((mul_34_17_n_8562 & mul_34_17_n_8230) | ((mul_34_17_n_8562 & mul_34_17_n_7667)
    | (mul_34_17_n_7667 & mul_34_17_n_8230)));
 assign mul_34_17_n_8984 = ((mul_34_17_n_8514 & mul_34_17_n_8409) | ((mul_34_17_n_8514 & mul_34_17_n_8030)
    | (mul_34_17_n_8030 & mul_34_17_n_8409)));
 assign mul_34_17_n_8982 = ((mul_34_17_n_8349 & mul_34_17_n_8419) | ((mul_34_17_n_8349 & mul_34_17_n_8378)
    | (mul_34_17_n_8378 & mul_34_17_n_8419)));
 assign mul_34_17_n_8950 = ~mul_34_17_n_8892;
 assign mul_34_17_n_8947 = ~mul_34_17_n_8946;
 assign mul_34_17_n_8945 = ~mul_34_17_n_8944;
 assign mul_34_17_n_8924 = ~mul_34_17_n_8925;
 assign mul_34_17_n_8920 = ~mul_34_17_n_8919;
 assign mul_34_17_n_8917 = ~mul_34_17_n_8916;
 assign mul_34_17_n_8912 = ~(mul_34_17_n_8592 | mul_34_17_n_8604);
 assign mul_34_17_n_8953 = ~(mul_34_17_n_8592 & mul_34_17_n_8604);
 assign mul_34_17_n_8911 = ~(mul_34_17_n_8643 & mul_34_17_n_8326);
 assign mul_34_17_n_8910 = ~(mul_34_17_n_8643 | mul_34_17_n_8326);
 assign mul_34_17_n_8909 = ~(mul_34_17_n_8602 & mul_34_17_n_8636);
 assign mul_34_17_n_8908 = ~(mul_34_17_n_8586 | mul_34_17_n_7626);
 assign mul_34_17_n_8907 = ~(mul_34_17_n_8616 | mul_34_17_n_8249);
 assign mul_34_17_n_8906 = ~(mul_34_17_n_8615 | mul_34_17_n_8250);
 assign mul_34_17_n_8905 = ~(mul_34_17_n_8706 | mul_34_17_n_8219);
 assign mul_34_17_n_8904 = ~(mul_34_17_n_364 | mul_34_17_n_8205);
 assign mul_34_17_n_8903 = ~(mul_34_17_n_363 | mul_34_17_n_7611);
 assign mul_34_17_n_8902 = ~(mul_34_17_n_8622 & mul_34_17_n_8673);
 assign mul_34_17_n_8901 = ~(mul_34_17_n_8489 ^ mul_34_17_n_7979);
 assign mul_34_17_n_8898 = ~((mul_34_17_n_7998 | mul_34_17_n_8202) & (mul_34_17_n_233 | mul_34_17_n_261));
 assign mul_34_17_n_8897 = (mul_34_17_n_8337 ^ mul_34_17_n_8380);
 assign mul_34_17_n_8952 = (mul_34_17_n_8030 ^ mul_34_17_n_8514);
 assign mul_34_17_n_8896 = ((mul_34_17_n_7902 | mul_34_17_n_7751) & (mul_34_17_n_8307 | mul_34_17_n_8452));
 assign mul_34_17_n_8895 = ~(mul_34_17_n_11380 ^ mul_34_17_n_11384);
 assign mul_34_17_n_8894 = ~(mul_34_17_n_8573 ^ mul_34_17_n_8269);
 assign mul_34_17_n_8893 = (mul_34_17_n_8348 ^ mul_34_17_n_8268);
 assign mul_34_17_n_8892 = ~(mul_34_17_n_8689 | mul_34_17_n_8274);
 assign mul_34_17_n_8891 = (mul_34_17_n_11376 ^ mul_34_17_n_11454);
 assign mul_34_17_n_8890 = ~(mul_34_17_n_8572 ^ mul_34_17_n_7915);
 assign mul_34_17_n_8889 = ~(mul_34_17_n_8301 ^ mul_34_17_n_7602);
 assign mul_34_17_n_8888 = (mul_34_17_n_8531 ^ mul_34_17_n_8403);
 assign mul_34_17_n_8887 = (mul_34_17_n_8355 ^ mul_34_17_n_8499);
 assign mul_34_17_n_8886 = ~(mul_34_17_n_8338 ^ mul_34_17_n_8509);
 assign mul_34_17_n_8885 = (mul_34_17_n_8349 ^ mul_34_17_n_8378);
 assign mul_34_17_n_8884 = (mul_34_17_n_8542 ^ mul_34_17_n_8523);
 assign mul_34_17_n_8883 = (mul_34_17_n_8032 ^ mul_34_17_n_8545);
 assign mul_34_17_n_8882 = (mul_34_17_n_231 ^ mul_34_17_n_8534);
 assign mul_34_17_n_8949 = ~(mul_34_17_n_8442 ^ mul_34_17_n_8151);
 assign mul_34_17_n_8948 = ~(mul_34_17_n_8447 ^ mul_34_17_n_7692);
 assign mul_34_17_n_8946 = ~(mul_34_17_n_8689 & mul_34_17_n_8274);
 assign mul_34_17_n_8944 = ~(mul_34_17_n_8433 ^ mul_34_17_n_7896);
 assign mul_34_17_n_8943 = ((mul_34_17_n_8235 & mul_34_17_n_7922) | ((mul_34_17_n_8235 & mul_34_17_n_8234)
    | (mul_34_17_n_8234 & mul_34_17_n_7922)));
 assign mul_34_17_n_8942 = ~((mul_34_17_n_8429 & ~mul_34_17_n_8421) | (mul_34_17_n_8574 & mul_34_17_n_8421));
 assign mul_34_17_n_8941 = ((mul_34_17_n_374 & mul_34_17_n_7769) | (mul_34_17_n_8480 & mul_34_17_n_7278));
 assign mul_34_17_n_8940 = ((mul_34_17_n_7887 & mul_34_17_n_247) | ((mul_34_17_n_7887 & mul_34_17_n_7885)
    | (mul_34_17_n_7885 & mul_34_17_n_247)));
 assign mul_34_17_n_8939 = ((mul_34_17_n_8141 & mul_34_17_n_7945) | ((mul_34_17_n_8141 & mul_34_17_n_7762)
    | (mul_34_17_n_7762 & mul_34_17_n_7945)));
 assign mul_34_17_n_8938 = ~(mul_34_17_n_8446 ^ mul_34_17_n_8142);
 assign mul_34_17_n_8937 = ((mul_34_17_n_8209 & mul_34_17_n_8071) | (mul_34_17_n_8478 & mul_34_17_n_7646));
 assign mul_34_17_n_8936 = ((mul_34_17_n_7998 & mul_34_17_n_233) | ((mul_34_17_n_7998 & mul_34_17_n_8253)
    | (mul_34_17_n_8253 & mul_34_17_n_233)));
 assign mul_34_17_n_8935 = ((mul_34_17_n_8277 & mul_34_17_n_8258) | ((mul_34_17_n_8277 & mul_34_17_n_7801)
    | (mul_34_17_n_7801 & mul_34_17_n_8258)));
 assign mul_34_17_n_8934 = ~(mul_34_17_n_8465 | (mul_34_17_n_8466 | (mul_34_17_n_8207 | mul_34_17_n_7970)));
 assign mul_34_17_n_8933 = ~((mul_34_17_n_368 & mul_34_17_n_8066) | (mul_34_17_n_8464 & mul_34_17_n_7607));
 assign mul_34_17_n_8932 = ~(mul_34_17_n_253 ^ mul_34_17_n_7734);
 assign mul_34_17_n_8931 = ((mul_34_17_n_7865 & mul_34_17_n_11420) | ((mul_34_17_n_7865 & mul_34_17_n_8255)
    | (mul_34_17_n_8255 & mul_34_17_n_11420)));
 assign mul_34_17_n_8930 = ~(mul_34_17_n_8441 ^ mul_34_17_n_7457);
 assign mul_34_17_n_8929 = ~(mul_34_17_n_8435 ^ mul_34_17_n_8340);
 assign mul_34_17_n_8928 = ((mul_34_17_n_8233 & mul_34_17_n_8555) | ((mul_34_17_n_8233 & mul_34_17_n_7752)
    | (mul_34_17_n_7752 & mul_34_17_n_8555)));
 assign mul_34_17_n_8927 = ~(mul_34_17_n_8439 ^ mul_34_17_n_8238);
 assign mul_34_17_n_8926 = ((mul_34_17_n_8022 & mul_34_17_n_8050) | ((mul_34_17_n_8022 & mul_34_17_n_8239)
    | (mul_34_17_n_8239 & mul_34_17_n_8050)));
 assign mul_34_17_n_8925 = ~(mul_34_17_n_8288 ^ mul_34_17_n_7764);
 assign mul_34_17_n_8923 = ((mul_34_17_n_8120 & mul_34_17_n_7558) | (mul_34_17_n_8475 & mul_34_17_n_7261));
 assign mul_34_17_n_8922 = ~(mul_34_17_n_8293 ^ mul_34_17_n_8136);
 assign mul_34_17_n_8921 = (mul_34_17_n_8552 ^ mul_34_17_n_8496);
 assign mul_34_17_n_8919 = ((mul_34_17_n_8010 & mul_34_17_n_8565) | ((mul_34_17_n_8010 & mul_34_17_n_8040)
    | (mul_34_17_n_8040 & mul_34_17_n_8565)));
 assign mul_34_17_n_8918 = ((mul_34_17_n_380 & mul_34_17_n_8056) | (mul_34_17_n_8479 & mul_34_17_n_7651));
 assign mul_34_17_n_8916 = ~(mul_34_17_n_8444 ^ mul_34_17_n_8004);
 assign mul_34_17_n_8915 = (mul_34_17_n_8571 ^ mul_34_17_n_7745);
 assign mul_34_17_n_8914 = (mul_34_17_n_8570 ^ mul_34_17_n_8261);
 assign mul_34_17_n_8913 = ~(mul_34_17_n_8434 ^ mul_34_17_n_8270);
 assign mul_34_17_n_8859 = ~mul_34_17_n_11342;
 assign mul_34_17_n_8856 = ~mul_34_17_n_259;
 assign mul_34_17_n_8847 = ~mul_34_17_n_8846;
 assign mul_34_17_n_8840 = ~mul_34_17_n_8839;
 assign mul_34_17_n_8831 = ~mul_34_17_n_8830;
 assign mul_34_17_n_8828 = ~mul_34_17_n_266;
 assign mul_34_17_n_8827 = ~mul_34_17_n_8826;
 assign mul_34_17_n_8825 = ~(mul_34_17_n_8330 ^ mul_34_17_n_8329);
 assign mul_34_17_n_8824 = ~(mul_34_17_n_8341 ^ mul_34_17_n_8013);
 assign mul_34_17_n_8823 = (mul_34_17_n_8411 ^ mul_34_17_n_8372);
 assign mul_34_17_n_8822 = ~((mul_34_17_n_6902 & (~mul_34_17_n_7895 & ~mul_34_17_n_8178)) | ((mul_34_17_n_6903
    & (mul_34_17_n_7895 & ~mul_34_17_n_8178)) | (mul_34_17_n_8449 & mul_34_17_n_8178)));
 assign mul_34_17_n_8821 = (mul_34_17_n_8158 ^ mul_34_17_n_8377);
 assign mul_34_17_n_8820 = (mul_34_17_n_8519 ^ mul_34_17_n_227);
 assign mul_34_17_n_8819 = (mul_34_17_n_8527 ^ mul_34_17_n_8388);
 assign mul_34_17_n_8818 = (mul_34_17_n_8541 ^ mul_34_17_n_7860);
 assign mul_34_17_n_8817 = (mul_34_17_n_8357 ^ mul_34_17_n_8358);
 assign mul_34_17_n_8816 = (mul_34_17_n_11370 ^ mul_34_17_n_8343);
 assign mul_34_17_n_8815 = (mul_34_17_n_8506 ^ mul_34_17_n_8554);
 assign mul_34_17_n_8814 = (mul_34_17_n_8360 ^ mul_34_17_n_8408);
 assign mul_34_17_n_8813 = (mul_34_17_n_8398 ^ mul_34_17_n_11625);
 assign mul_34_17_n_8881 = ~(mul_34_17_n_8367 ^ mul_34_17_n_7427);
 assign mul_34_17_n_8812 = (mul_34_17_n_8368 ^ mul_34_17_n_8009);
 assign mul_34_17_n_8880 = (mul_34_17_n_8384 ^ mul_34_17_n_8415);
 assign mul_34_17_n_8811 = ~(mul_34_17_n_8399 ^ mul_34_17_n_7877);
 assign mul_34_17_n_8810 = (mul_34_17_n_8418 ^ mul_34_17_n_7899);
 assign mul_34_17_n_8809 = (mul_34_17_n_8420 ^ mul_34_17_n_8354);
 assign mul_34_17_n_8808 = ~(mul_34_17_n_8564 ^ mul_34_17_n_8392);
 assign mul_34_17_n_8879 = ~(mul_34_17_n_8292 ^ mul_34_17_n_7583);
 assign mul_34_17_n_8807 = (mul_34_17_n_8364 ^ mul_34_17_n_8263);
 assign mul_34_17_n_8878 = ~(mul_34_17_n_8305 ^ mul_34_17_n_8143);
 assign mul_34_17_n_8806 = (mul_34_17_n_8342 ^ mul_34_17_n_8259);
 assign mul_34_17_n_8877 = ((mul_34_17_n_8113 & mul_34_17_n_7923) | (mul_34_17_n_8472 & mul_34_17_n_7635));
 assign mul_34_17_n_8876 = ~(mul_34_17_n_8303 ^ mul_34_17_n_7471);
 assign mul_34_17_n_8875 = ~((mul_34_17_n_7416 & (~mul_34_17_n_7855 & ~mul_34_17_n_7497)) | ((mul_34_17_n_7415
    & (mul_34_17_n_7855 & ~mul_34_17_n_7497)) | (mul_34_17_n_8313 & mul_34_17_n_7497)));
 assign mul_34_17_n_8874 = ~(mul_34_17_n_8300 ^ mul_34_17_n_7551);
 assign mul_34_17_n_8873 = ~(mul_34_17_n_8284 ^ mul_34_17_n_7318);
 assign mul_34_17_n_8872 = ~(mul_34_17_n_8255 ^ mul_34_17_n_8289);
 assign mul_34_17_n_8870 = ~(mul_34_17_n_8290 ^ mul_34_17_n_7888);
 assign mul_34_17_n_8869 = ((mul_34_17_n_8012 & mul_34_17_n_11424) | ((mul_34_17_n_8012 & mul_34_17_n_8143)
    | (mul_34_17_n_8143 & mul_34_17_n_11424)));
 assign mul_34_17_n_8805 = ~(mul_34_17_n_8424 ^ mul_34_17_n_7890);
 assign mul_34_17_n_8868 = ~(mul_34_17_n_8302 ^ mul_34_17_n_7757);
 assign mul_34_17_n_8867 = ~((mul_34_17_n_367 & mul_34_17_n_7929) | (mul_34_17_n_8473 & mul_34_17_n_7639));
 assign mul_34_17_n_8866 = ~(mul_34_17_n_8294 ^ mul_34_17_n_8156);
 assign mul_34_17_n_8865 = ~(mul_34_17_n_8396 ^ mul_34_17_n_7681);
 assign mul_34_17_n_8864 = ~((mul_34_17_n_218 & (~mul_34_17_n_11470 & ~mul_34_17_n_7728)) | ((mul_34_17_n_7993
    & (mul_34_17_n_11470 & ~mul_34_17_n_7728)) | (mul_34_17_n_8450 & mul_34_17_n_7728)));
 assign mul_34_17_n_8863 = ~((mul_34_17_n_5512 & (~mul_34_17_n_6912 & ~mul_34_17_n_8436)) | ((mul_34_17_n_5513
    & (mul_34_17_n_6912 & ~mul_34_17_n_8436)) | (mul_34_17_n_7773 & mul_34_17_n_8436)));
 assign mul_34_17_n_8860 = ~((mul_34_17_n_7835 & (~mul_34_17_n_7843 & ~mul_34_17_n_7474)) | ((mul_34_17_n_7834
    & (mul_34_17_n_7843 & ~mul_34_17_n_7474)) | (mul_34_17_n_8458 & mul_34_17_n_7474)));
 assign mul_34_17_n_8855 = ((mul_34_17_n_378 & mul_34_17_n_7937) | (mul_34_17_n_8467 & mul_34_17_n_7621));
 assign mul_34_17_n_8854 = ((mul_34_17_n_11635 & mul_34_17_n_11430) | ((mul_34_17_n_11635 & mul_34_17_n_8136)
    | (mul_34_17_n_8136 & mul_34_17_n_11430)));
 assign mul_34_17_n_8853 = ~(mul_34_17_n_8304 ^ mul_34_17_n_8020);
 assign mul_34_17_n_8852 = ~(mul_34_17_n_8299 ^ mul_34_17_n_8059);
 assign mul_34_17_n_8851 = ~((mul_34_17_n_8115 & mul_34_17_n_7943) | (mul_34_17_n_8321 & mul_34_17_n_7609));
 assign mul_34_17_n_8850 = ~(mul_34_17_n_8407 ^ mul_34_17_n_8008);
 assign mul_34_17_n_8849 = ~(mul_34_17_n_8286 ^ mul_34_17_n_8374);
 assign mul_34_17_n_8848 = (mul_34_17_n_8383 ^ mul_34_17_n_8266);
 assign mul_34_17_n_8846 = ((mul_34_17_n_11631 & mul_34_17_n_11627) | ((mul_34_17_n_11631 & mul_34_17_n_8142)
    | (mul_34_17_n_8142 & mul_34_17_n_11627)));
 assign mul_34_17_n_8845 = ~(mul_34_17_n_7894 ^ mul_34_17_n_8291);
 assign mul_34_17_n_8844 = (mul_34_17_n_8371 ^ mul_34_17_n_8416);
 assign mul_34_17_n_8843 = ((mul_34_17_n_8126 & mul_34_17_n_8131) | ((mul_34_17_n_8126 & mul_34_17_n_7927)
    | (mul_34_17_n_7927 & mul_34_17_n_8131)));
 assign mul_34_17_n_8842 = ~(mul_34_17_n_8426 ^ mul_34_17_n_7535);
 assign mul_34_17_n_8841 = ~(mul_34_17_n_8296 ^ mul_34_17_n_7702);
 assign mul_34_17_n_8839 = (mul_34_17_n_8427 ^ mul_34_17_n_7858);
 assign mul_34_17_n_8838 = ~(mul_34_17_n_8297 ^ mul_34_17_n_8265);
 assign mul_34_17_n_8835 = ((mul_34_17_n_372 & mul_34_17_n_7924) | (mul_34_17_n_8474 & mul_34_17_n_7610));
 assign mul_34_17_n_8834 = ~((mul_34_17_n_219 & ~mul_34_17_n_160) | (mul_34_17_n_8453 & mul_34_17_n_160));
 assign mul_34_17_n_8830 = ((mul_34_17_n_11444 & mul_34_17_n_8567) | ((mul_34_17_n_11444 & mul_34_17_n_8144)
    | (mul_34_17_n_8144 & mul_34_17_n_8567)));
 assign mul_34_17_n_8829 = ((mul_34_17_n_8246 & mul_34_17_n_8399) | ((mul_34_17_n_8246 & mul_34_17_n_7878)
    | (mul_34_17_n_7878 & mul_34_17_n_8399)));
 assign mul_34_17_n_8826 = ((mul_34_17_n_7872 & mul_34_17_n_8412) | ((mul_34_17_n_7872 & mul_34_17_n_7876)
    | (mul_34_17_n_7876 & mul_34_17_n_8412)));
 assign mul_34_17_n_8799 = ~mul_34_17_n_8798;
 assign mul_34_17_n_8793 = ~mul_34_17_n_8792;
 assign mul_34_17_n_8791 = ~mul_34_17_n_8790;
 assign mul_34_17_n_8788 = ~mul_34_17_n_8787;
 assign mul_34_17_n_8785 = ~mul_34_17_n_8784;
 assign mul_34_17_n_8769 = ~mul_34_17_n_8768;
 assign mul_34_17_n_8765 = ~mul_34_17_n_8764;
 assign mul_34_17_n_8760 = ~mul_34_17_n_8761;
 assign mul_34_17_n_8754 = ~mul_34_17_n_251;
 assign mul_34_17_n_8742 = ~mul_34_17_n_8741;
 assign mul_34_17_n_8736 = ~mul_34_17_n_8735;
 assign mul_34_17_n_8728 = ~mul_34_17_n_8727;
 assign mul_34_17_n_8722 = ~mul_34_17_n_8721;
 assign mul_34_17_n_8719 = ~mul_34_17_n_8720;
 assign mul_34_17_n_8717 = ~(mul_34_17_n_8548 | mul_34_17_n_8226);
 assign mul_34_17_n_8716 = ~(mul_34_17_n_8548 & mul_34_17_n_8226);
 assign mul_34_17_n_8715 = ~(mul_34_17_n_371 | mul_34_17_n_7658);
 assign mul_34_17_n_8714 = ((mul_34_17_n_7842 | mul_34_17_n_7996) & (mul_34_17_n_8214 | mul_34_17_n_8215));
 assign mul_34_17_n_8713 = ~(mul_34_17_n_8468 | mul_34_17_n_7653);
 assign mul_34_17_n_8712 = ~(mul_34_17_n_370 | mul_34_17_n_7649);
 assign mul_34_17_n_8711 = ~(mul_34_17_n_228 ^ mul_34_17_n_8231);
 assign mul_34_17_n_8710 = ~(mul_34_17_n_8311 | mul_34_17_n_7633);
 assign mul_34_17_n_8709 = ~(mul_34_17_n_247 & mul_34_17_n_8429);
 assign mul_34_17_n_8708 = ~(mul_34_17_n_247 & mul_34_17_n_8187);
 assign mul_34_17_n_8707 = (mul_34_17_n_228 ^ mul_34_17_n_8231);
 assign mul_34_17_n_8706 = (mul_34_17_n_8229 ^ mul_34_17_n_7667);
 assign mul_34_17_n_8705 = ~(mul_34_17_n_366 | mul_34_17_n_7616);
 assign mul_34_17_n_8704 = ~(mul_34_17_n_365 | mul_34_17_n_7614);
 assign mul_34_17_n_8703 = ~(mul_34_17_n_8165 ^ mul_34_17_n_8070);
 assign mul_34_17_n_8701 = ~(mul_34_17_n_8230 ^ mul_34_17_n_7667);
 assign mul_34_17_n_8700 = ~(mul_34_17_n_8482 | mul_34_17_n_7664);
 assign mul_34_17_n_8699 = ((mul_34_17_n_6408 & mul_34_17_n_8279) | ((mul_34_17_n_6408 & mul_34_17_n_6687)
    | (mul_34_17_n_6687 & mul_34_17_n_8279)));
 assign mul_34_17_n_8698 = ~(mul_34_17_n_8421 & mul_34_17_n_8574);
 assign mul_34_17_n_8696 = (mul_34_17_n_8245 ^ mul_34_17_n_8062);
 assign mul_34_17_n_8804 = ((mul_34_17_n_7880 & mul_34_17_n_7583) | ((mul_34_17_n_7880 & mul_34_17_n_7756)
    | (mul_34_17_n_7756 & mul_34_17_n_7583)));
 assign mul_34_17_n_8803 = ~(mul_34_17_n_8134 ^ mul_34_17_n_7435);
 assign mul_34_17_n_8802 = ~(mul_34_17_n_8195 ^ mul_34_17_n_8154);
 assign mul_34_17_n_8801 = ~(mul_34_17_n_7489 ^ (mul_34_17_n_7794 ^ (mul_34_17_n_6804 ^ mul_34_17_n_5906)));
 assign mul_34_17_n_8695 = (mul_34_17_n_8233 ^ mul_34_17_n_7752);
 assign mul_34_17_n_8798 = ~(mul_34_17_n_8208 | (mul_34_17_n_7973 | (mul_34_17_n_8222 | mul_34_17_n_7601)));
 assign mul_34_17_n_8694 = (mul_34_17_n_8277 ^ mul_34_17_n_7801);
 assign mul_34_17_n_8693 = ~(mul_34_17_n_8490 | mul_34_17_n_7979);
 assign mul_34_17_n_8797 = ~(mul_34_17_n_8191 ^ mul_34_17_n_7317);
 assign mul_34_17_n_8692 = ((mul_34_17_n_11442 & mul_34_17_n_8271) | ((mul_34_17_n_11442 & mul_34_17_n_11440)
    | (mul_34_17_n_11440 & mul_34_17_n_8271)));
 assign mul_34_17_n_8796 = ((mul_34_17_n_8025 & mul_34_17_n_8264) | ((mul_34_17_n_8025 & mul_34_17_n_7759)
    | (mul_34_17_n_7759 & mul_34_17_n_8264)));
 assign mul_34_17_n_8795 = ((mul_34_17_n_7987 & mul_34_17_n_8228) | ((mul_34_17_n_7987 & mul_34_17_n_7716)
    | (mul_34_17_n_7716 & mul_34_17_n_8228)));
 assign mul_34_17_n_8794 = ~(mul_34_17_n_8180 ^ mul_34_17_n_7123);
 assign mul_34_17_n_8691 = (mul_34_17_n_8235 ^ mul_34_17_n_7922);
 assign mul_34_17_n_8792 = ((mul_34_17_n_7938 & mul_34_17_n_7156) | (mul_34_17_n_8272 & mul_34_17_n_8188));
 assign mul_34_17_n_8790 = ((mul_34_17_n_8007 & mul_34_17_n_8153) | ((mul_34_17_n_8007 & mul_34_17_n_8028)
    | (mul_34_17_n_8028 & mul_34_17_n_8153)));
 assign mul_34_17_n_8789 = ((mul_34_17_n_8053 & mul_34_17_n_11410) | ((mul_34_17_n_8053 & mul_34_17_n_11418)
    | (mul_34_17_n_11418 & mul_34_17_n_11410)));
 assign mul_34_17_n_8787 = ((mul_34_17_n_7839 & mul_34_17_n_7846) | ((mul_34_17_n_7839 & mul_34_17_n_8049)
    | (mul_34_17_n_8049 & mul_34_17_n_7846)));
 assign mul_34_17_n_8786 = ((mul_34_17_n_182 & mul_34_17_n_11629) | ((mul_34_17_n_182 & mul_34_17_n_8003)
    | (mul_34_17_n_8003 & mul_34_17_n_11629)));
 assign mul_34_17_n_8784 = ~(mul_34_17_n_8179 ^ mul_34_17_n_7748);
 assign mul_34_17_n_8783 = ((mul_34_17_n_7897 & mul_34_17_n_8048) | ((mul_34_17_n_7897 & mul_34_17_n_7719)
    | (mul_34_17_n_7719 & mul_34_17_n_8048)));
 assign mul_34_17_n_8782 = ~(mul_34_17_n_8189 ^ mul_34_17_n_7697);
 assign mul_34_17_n_8780 = ((mul_34_17_n_7986 & mul_34_17_n_11466) | ((mul_34_17_n_7986 & mul_34_17_n_7492)
    | (mul_34_17_n_7492 & mul_34_17_n_11466)));
 assign mul_34_17_n_8779 = ((mul_34_17_n_7875 & mul_34_17_n_223) | ((mul_34_17_n_7875 & mul_34_17_n_7744)
    | (mul_34_17_n_7744 & mul_34_17_n_223)));
 assign mul_34_17_n_8777 = ~(mul_34_17_n_8182 ^ mul_34_17_n_7717);
 assign mul_34_17_n_8776 = ((mul_34_17_n_7594 & mul_34_17_n_8155) | ((mul_34_17_n_7594 & mul_34_17_n_7797)
    | (mul_34_17_n_7797 & mul_34_17_n_8155)));
 assign mul_34_17_n_8775 = ((mul_34_17_n_8002 & mul_34_17_n_8065) | ((mul_34_17_n_8002 & mul_34_17_n_7743)
    | (mul_34_17_n_7743 & mul_34_17_n_8065)));
 assign mul_34_17_n_8773 = ~(mul_34_17_n_8095 ^ mul_34_17_n_7576);
 assign mul_34_17_n_8771 = ~(mul_34_17_n_8183 ^ mul_34_17_n_7783);
 assign mul_34_17_n_8770 = ~(mul_34_17_n_8276 ^ mul_34_17_n_7788);
 assign mul_34_17_n_8768 = ((mul_34_17_n_11478 & mul_34_17_n_11464) | ((mul_34_17_n_11478 & mul_34_17_n_7701)
    | (mul_34_17_n_7701 & mul_34_17_n_11464)));
 assign mul_34_17_n_8767 = (mul_34_17_n_8256 ^ mul_34_17_n_7898);
 assign mul_34_17_n_8766 = ~((mul_34_17_n_7703 & mul_34_17_n_155) | (mul_34_17_n_8200 & mul_34_17_n_7276));
 assign mul_34_17_n_8764 = ((mul_34_17_n_7983 & mul_34_17_n_215) | ((mul_34_17_n_7983 & mul_34_17_n_160)
    | (mul_34_17_n_160 & mul_34_17_n_215)));
 assign mul_34_17_n_8763 = ((mul_34_17_n_8031 & mul_34_17_n_8044) | ((mul_34_17_n_8031 & mul_34_17_n_7692)
    | (mul_34_17_n_7692 & mul_34_17_n_8044)));
 assign mul_34_17_n_8762 = ~(mul_34_17_n_8190 ^ mul_34_17_n_11633);
 assign mul_34_17_n_8761 = ~(mul_34_17_n_8275 ^ mul_34_17_n_7767);
 assign mul_34_17_n_8759 = ~(mul_34_17_n_8176 ^ mul_34_17_n_7363);
 assign mul_34_17_n_8758 = ((mul_34_17_n_7993 & mul_34_17_n_11470) | ((mul_34_17_n_7993 & mul_34_17_n_7729)
    | (mul_34_17_n_7729 & mul_34_17_n_11470)));
 assign mul_34_17_n_8757 = ~(mul_34_17_n_8192 ^ mul_34_17_n_7795);
 assign mul_34_17_n_8756 = ((mul_34_17_n_8055 & mul_34_17_n_7852) | ((mul_34_17_n_8055 & mul_34_17_n_7981)
    | (mul_34_17_n_7981 & mul_34_17_n_7852)));
 assign mul_34_17_n_8755 = ~(mul_34_17_n_8175 ^ mul_34_17_n_7731);
 assign mul_34_17_n_8753 = ((mul_34_17_n_384 & mul_34_17_n_7850) | ((mul_34_17_n_384 & mul_34_17_n_7838)
    | (mul_34_17_n_7838 & mul_34_17_n_7850)));
 assign mul_34_17_n_8752 = ((mul_34_17_n_11460 & mul_34_17_n_7908) | ((mul_34_17_n_11460 & mul_34_17_n_7894)
    | (mul_34_17_n_7894 & mul_34_17_n_7908)));
 assign mul_34_17_n_8751 = ~(mul_34_17_n_8174 ^ mul_34_17_n_7452);
 assign mul_34_17_n_8750 = ((mul_34_17_n_375 & mul_34_17_n_149) | (mul_34_17_n_8221 & mul_34_17_n_6451));
 assign mul_34_17_n_8749 = ~(mul_34_17_n_8196 ^ mul_34_17_n_11500);
 assign mul_34_17_n_8748 = ~(mul_34_17_n_8186 ^ mul_34_17_n_7137);
 assign mul_34_17_n_8747 = ~(mul_34_17_n_8089 ^ mul_34_17_n_7713);
 assign mul_34_17_n_8746 = ~(mul_34_17_n_8102 ^ mul_34_17_n_7462);
 assign mul_34_17_n_8745 = ((mul_34_17_n_11448 & mul_34_17_n_8151) | ((mul_34_17_n_11448 & mul_34_17_n_11392)
    | (mul_34_17_n_11392 & mul_34_17_n_8151)));
 assign mul_34_17_n_8744 = ((mul_34_17_n_165 & mul_34_17_n_8052) | ((mul_34_17_n_165 & mul_34_17_n_8005)
    | (mul_34_17_n_8005 & mul_34_17_n_8052)));
 assign mul_34_17_n_8743 = ~(mul_34_17_n_8073 ^ mul_34_17_n_7726);
 assign mul_34_17_n_8741 = ((mul_34_17_n_229 & mul_34_17_n_8265) | ((mul_34_17_n_229 & mul_34_17_n_11446)
    | (mul_34_17_n_11446 & mul_34_17_n_8265)));
 assign mul_34_17_n_8740 = ((mul_34_17_n_7864 & mul_34_17_n_7786) | ((mul_34_17_n_7864 & mul_34_17_n_7319)
    | (mul_34_17_n_7319 & mul_34_17_n_7786)));
 assign mul_34_17_n_8739 = ((mul_34_17_n_8123 & mul_34_17_n_8057) | (mul_34_17_n_8210 & mul_34_17_n_7959));
 assign mul_34_17_n_8738 = ((mul_34_17_n_11452 & mul_34_17_n_8156) | ((mul_34_17_n_11452 & mul_34_17_n_11450)
    | (mul_34_17_n_11450 & mul_34_17_n_8156)));
 assign mul_34_17_n_8737 = ((mul_34_17_n_11402 & mul_34_17_n_8261) | ((mul_34_17_n_11402 & mul_34_17_n_7685)
    | (mul_34_17_n_7685 & mul_34_17_n_8261)));
 assign mul_34_17_n_8735 = ((mul_34_17_n_11398 & mul_34_17_n_8267) | ((mul_34_17_n_11398 & mul_34_17_n_7538)
    | (mul_34_17_n_7538 & mul_34_17_n_8267)));
 assign mul_34_17_n_8734 = ((mul_34_17_n_11414 & mul_34_17_n_11404) | ((mul_34_17_n_11414 & mul_34_17_n_8019)
    | (mul_34_17_n_8019 & mul_34_17_n_11404)));
 assign mul_34_17_n_8733 = ~(mul_34_17_n_8092 ^ mul_34_17_n_7766);
 assign mul_34_17_n_8732 = ~((mul_34_17_n_8033 & mul_34_17_n_7755) | (mul_34_17_n_8217 & mul_34_17_n_8260));
 assign mul_34_17_n_8731 = ~(mul_34_17_n_8185 ^ mul_34_17_n_7573);
 assign mul_34_17_n_8730 = ~(mul_34_17_n_8090 ^ mul_34_17_n_7302);
 assign mul_34_17_n_8727 = (mul_34_17_n_8273 ^ mul_34_17_n_7739);
 assign mul_34_17_n_8726 = ((mul_34_17_n_8017 & mul_34_17_n_11426) | ((mul_34_17_n_8017 & mul_34_17_n_7757)
    | (mul_34_17_n_7757 & mul_34_17_n_11426)));
 assign mul_34_17_n_8724 = ((mul_34_17_n_11474 & mul_34_17_n_11468) | ((mul_34_17_n_11474 & mul_34_17_n_7700)
    | (mul_34_17_n_7700 & mul_34_17_n_11468)));
 assign mul_34_17_n_8723 = ((mul_34_17_n_8015 & mul_34_17_n_11428) | ((mul_34_17_n_8015 & mul_34_17_n_7536)
    | (mul_34_17_n_7536 & mul_34_17_n_11428)));
 assign mul_34_17_n_8721 = (mul_34_17_n_8278 ^ mul_34_17_n_7566);
 assign mul_34_17_n_8720 = ~(mul_34_17_n_8184 ^ mul_34_17_n_7330);
 assign mul_34_17_n_8676 = ~mul_34_17_n_8675;
 assign mul_34_17_n_8669 = ~mul_34_17_n_8668;
 assign mul_34_17_n_8660 = ~mul_34_17_n_256;
 assign mul_34_17_n_8656 = ~mul_34_17_n_8655;
 assign mul_34_17_n_8646 = ~mul_34_17_n_8647;
 assign mul_34_17_n_8643 = ~mul_34_17_n_8642;
 assign mul_34_17_n_8637 = ~mul_34_17_n_8636;
 assign mul_34_17_n_8635 = ~mul_34_17_n_11364;
 assign mul_34_17_n_8627 = ~mul_34_17_n_8628;
 assign mul_34_17_n_8623 = ~mul_34_17_n_8622;
 assign mul_34_17_n_8616 = ~mul_34_17_n_8615;
 assign mul_34_17_n_8608 = ~mul_34_17_n_8607;
 assign mul_34_17_n_8605 = ~mul_34_17_n_11368;
 assign mul_34_17_n_8603 = ~mul_34_17_n_8604;
 assign mul_34_17_n_8601 = ~mul_34_17_n_8602;
 assign mul_34_17_n_8600 = ~mul_34_17_n_8599;
 assign mul_34_17_n_8597 = ~mul_34_17_n_8596;
 assign mul_34_17_n_8594 = ~mul_34_17_n_8595;
 assign mul_34_17_n_8591 = ~mul_34_17_n_8592;
 assign mul_34_17_n_8590 = ~(mul_34_17_n_8228 ^ mul_34_17_n_164);
 assign mul_34_17_n_8589 = ~(mul_34_17_n_8130 ^ mul_34_17_n_180);
 assign mul_34_17_n_8587 = ~(mul_34_17_n_8126 ^ mul_34_17_n_8131);
 assign mul_34_17_n_8586 = ~(mul_34_17_n_8131 ^ mul_34_17_n_8126);
 assign mul_34_17_n_8585 = ~(mul_34_17_n_8129 ^ mul_34_17_n_7422);
 assign mul_34_17_n_8584 = (mul_34_17_n_8149 ^ mul_34_17_n_7712);
 assign mul_34_17_n_8583 = (mul_34_17_n_11444 ^ mul_34_17_n_8144);
 assign mul_34_17_n_8690 = (mul_34_17_n_11400 ^ mul_34_17_n_8262);
 assign mul_34_17_n_8689 = ~(mul_34_17_n_7373 ^ mul_34_17_n_8193);
 assign mul_34_17_n_8688 = ~(mul_34_17_n_8163 ^ mul_34_17_n_7918);
 assign mul_34_17_n_8687 = ~(mul_34_17_n_8083 ^ mul_34_17_n_7704);
 assign mul_34_17_n_8582 = (mul_34_17_n_8260 ^ mul_34_17_n_8033);
 assign mul_34_17_n_8581 = (mul_34_17_n_232 ^ mul_34_17_n_8157);
 assign mul_34_17_n_8580 = (mul_34_17_n_8145 ^ mul_34_17_n_11388);
 assign mul_34_17_n_8579 = ~(mul_34_17_n_8241 ^ mul_34_17_n_7906);
 assign mul_34_17_n_8686 = ((mul_34_17_n_7832 & mul_34_17_n_7853) | ((mul_34_17_n_7832 & mul_34_17_n_7483)
    | (mul_34_17_n_7483 & mul_34_17_n_7853)));
 assign mul_34_17_n_8578 = (mul_34_17_n_8170 ^ mul_34_17_n_7518);
 assign mul_34_17_n_8684 = ((mul_34_17_n_11416 & mul_34_17_n_7854) | ((mul_34_17_n_11416 & mul_34_17_n_7934)
    | (mul_34_17_n_7934 & mul_34_17_n_7854)));
 assign mul_34_17_n_8682 = ~(mul_34_17_n_8088 ^ mul_34_17_n_7905);
 assign mul_34_17_n_8680 = ((mul_34_17_n_11639 & mul_34_17_n_11422) | ((mul_34_17_n_11639 & mul_34_17_n_7764)
    | (mul_34_17_n_7764 & mul_34_17_n_11422)));
 assign mul_34_17_n_8678 = ~((mul_34_17_n_7675 & (~mul_34_17_n_7441 & ~mul_34_17_n_7493)) | ((mul_34_17_n_7674
    & (mul_34_17_n_7441 & ~mul_34_17_n_7493)) | (mul_34_17_n_8108 & mul_34_17_n_7493)));
 assign mul_34_17_n_8677 = ((mul_34_17_n_7805 & mul_34_17_n_7807) | ((mul_34_17_n_7805 & mul_34_17_n_7457)
    | (mul_34_17_n_7457 & mul_34_17_n_7807)));
 assign mul_34_17_n_8675 = ((mul_34_17_n_373 & mul_34_17_n_7593) | (mul_34_17_n_8118 & mul_34_17_n_7390));
 assign mul_34_17_n_8674 = ((mul_34_17_n_7836 & mul_34_17_n_8130) | ((mul_34_17_n_7836 & mul_34_17_n_7454)
    | (mul_34_17_n_7454 & mul_34_17_n_8130)));
 assign mul_34_17_n_8673 = ~(mul_34_17_n_8135 ^ mul_34_17_n_7423);
 assign mul_34_17_n_8672 = ((mul_34_17_n_377 & mul_34_17_n_7584) | (mul_34_17_n_8204 & mul_34_17_n_7248));
 assign mul_34_17_n_8671 = ~((mul_34_17_n_7673 & (~mul_34_17_n_167 & ~mul_34_17_n_7753)) | ((mul_34_17_n_7672
    & (mul_34_17_n_167 & ~mul_34_17_n_7753)) | (mul_34_17_n_8201 & mul_34_17_n_7753)));
 assign mul_34_17_n_8670 = ~(mul_34_17_n_8133 ^ mul_34_17_n_7424);
 assign mul_34_17_n_8668 = ~((mul_34_17_n_8218 & ~mul_34_17_n_8046) | (mul_34_17_n_8199 & mul_34_17_n_8046));
 assign mul_34_17_n_8666 = ((mul_34_17_n_11458 & mul_34_17_n_11432) | ((mul_34_17_n_11458 & mul_34_17_n_7551)
    | (mul_34_17_n_7551 & mul_34_17_n_11432)));
 assign mul_34_17_n_8664 = ((mul_34_17_n_8057 & mul_34_17_n_7684) | ((mul_34_17_n_8057 & mul_34_17_n_7414)
    | (mul_34_17_n_7414 & mul_34_17_n_7684)));
 assign mul_34_17_n_8663 = ((mul_34_17_n_7925 & mul_34_17_n_7429) | ((mul_34_17_n_7925 & mul_34_17_n_7411)
    | (mul_34_17_n_7411 & mul_34_17_n_7429)));
 assign mul_34_17_n_8662 = ~(mul_34_17_n_8082 ^ mul_34_17_n_7555);
 assign mul_34_17_n_8661 = ~(mul_34_17_n_8096 ^ mul_34_17_n_7315);
 assign mul_34_17_n_8659 = ((mul_34_17_n_7882 & mul_34_17_n_8148) | ((mul_34_17_n_7882 & mul_34_17_n_7869)
    | (mul_34_17_n_7869 & mul_34_17_n_8148)));
 assign mul_34_17_n_8658 = ~(mul_34_17_n_8086 ^ mul_34_17_n_11498);
 assign mul_34_17_n_8657 = ((mul_34_17_n_11462 & mul_34_17_n_8059) | ((mul_34_17_n_11462 & mul_34_17_n_11390)
    | (mul_34_17_n_11390 & mul_34_17_n_8059)));
 assign mul_34_17_n_8655 = ~(mul_34_17_n_8060 ^ mul_34_17_n_8166);
 assign mul_34_17_n_8654 = ~(mul_34_17_n_8106 ^ mul_34_17_n_7556);
 assign mul_34_17_n_8653 = (mul_34_17_n_8172 ^ mul_34_17_n_202);
 assign mul_34_17_n_8652 = ~(mul_34_17_n_8105 ^ mul_34_17_n_7705);
 assign mul_34_17_n_8651 = (mul_34_17_n_8173 ^ mul_34_17_n_7085);
 assign mul_34_17_n_8650 = ((mul_34_17_n_7857 & mul_34_17_n_11436) | ((mul_34_17_n_7857 & mul_34_17_n_163)
    | (mul_34_17_n_163 & mul_34_17_n_11436)));
 assign mul_34_17_n_8649 = ~(mul_34_17_n_7336 ^ mul_34_17_n_8103);
 assign mul_34_17_n_8648 = ~(mul_34_17_n_8080 ^ mul_34_17_n_7097);
 assign mul_34_17_n_8647 = (mul_34_17_n_7066 ^ mul_34_17_n_8171);
 assign mul_34_17_n_8645 = ~(mul_34_17_n_8098 ^ mul_34_17_n_7490);
 assign mul_34_17_n_8644 = ((mul_34_17_n_7933 & mul_34_17_n_11408) | ((mul_34_17_n_7933 & mul_34_17_n_11412)
    | (mul_34_17_n_11412 & mul_34_17_n_11408)));
 assign mul_34_17_n_8642 = ~(mul_34_17_n_8152 ^ mul_34_17_n_8236);
 assign mul_34_17_n_8641 = ((mul_34_17_n_11479 & mul_34_17_n_11406) | ((mul_34_17_n_11479 & mul_34_17_n_7900)
    | (mul_34_17_n_7900 & mul_34_17_n_11406)));
 assign mul_34_17_n_8640 = ((mul_34_17_n_11396 & mul_34_17_n_11438) | ((mul_34_17_n_11396 & mul_34_17_n_7535)
    | (mul_34_17_n_7535 & mul_34_17_n_11438)));
 assign mul_34_17_n_8639 = ~(mul_34_17_n_8078 ^ mul_34_17_n_7091);
 assign mul_34_17_n_8638 = ~(mul_34_17_n_8077 ^ mul_34_17_n_7087);
 assign mul_34_17_n_8636 = ~(mul_34_17_n_8181 ^ mul_34_17_n_7068);
 assign mul_34_17_n_8633 = ((mul_34_17_n_8016 & mul_34_17_n_7911) | ((mul_34_17_n_8016 & mul_34_17_n_7541)
    | (mul_34_17_n_7541 & mul_34_17_n_7911)));
 assign mul_34_17_n_8577 = (mul_34_17_n_8160 ^ mul_34_17_n_8161);
 assign mul_34_17_n_8632 = ~(mul_34_17_n_8074 ^ mul_34_17_n_7585);
 assign mul_34_17_n_8631 = ((mul_34_17_n_11476 & mul_34_17_n_11472) | ((mul_34_17_n_11476 & mul_34_17_n_159)
    | (mul_34_17_n_159 & mul_34_17_n_11472)));
 assign mul_34_17_n_8630 = ~(mul_34_17_n_8094 ^ mul_34_17_n_7309);
 assign mul_34_17_n_8629 = ((mul_34_17_n_7929 & mul_34_17_n_11489) | ((mul_34_17_n_7929 & mul_34_17_n_7410)
    | (mul_34_17_n_7410 & mul_34_17_n_11489)));
 assign mul_34_17_n_8628 = ~(mul_34_17_n_8159 ^ mul_34_17_n_7592);
 assign mul_34_17_n_8626 = ~(mul_34_17_n_8167 ^ mul_34_17_n_11637);
 assign mul_34_17_n_8625 = ((mul_34_17_n_11481 & mul_34_17_n_8224) | ((mul_34_17_n_11481 & mul_34_17_n_224)
    | (mul_34_17_n_224 & mul_34_17_n_8224)));
 assign mul_34_17_n_8624 = ~(mul_34_17_n_8081 ^ mul_34_17_n_7339);
 assign mul_34_17_n_8622 = ~(mul_34_17_n_8076 ^ mul_34_17_n_7465);
 assign mul_34_17_n_8621 = ((mul_34_17_n_7871 & mul_34_17_n_7680) | ((mul_34_17_n_7871 & mul_34_17_n_7119)
    | (mul_34_17_n_7119 & mul_34_17_n_7680)));
 assign mul_34_17_n_8620 = ~(mul_34_17_n_8093 ^ mul_34_17_n_7378);
 assign mul_34_17_n_8619 = ((mul_34_17_n_8024 & mul_34_17_n_11434) | ((mul_34_17_n_8024 & mul_34_17_n_8021)
    | (mul_34_17_n_8021 & mul_34_17_n_11434)));
 assign mul_34_17_n_8618 = ((mul_34_17_n_7884 & mul_34_17_n_7903) | ((mul_34_17_n_7884 & mul_34_17_n_7888)
    | (mul_34_17_n_7888 & mul_34_17_n_7903)));
 assign mul_34_17_n_8617 = ~(mul_34_17_n_8099 ^ mul_34_17_n_7129);
 assign mul_34_17_n_8615 = ~(mul_34_17_n_8162 ^ mul_34_17_n_7781);
 assign mul_34_17_n_8576 = ~(mul_34_17_n_8168 ^ mul_34_17_n_7567);
 assign mul_34_17_n_8613 = ~(mul_34_17_n_8085 ^ mul_34_17_n_7128);
 assign mul_34_17_n_8575 = (mul_34_17_n_8169 ^ mul_34_17_n_7515);
 assign mul_34_17_n_8612 = ((mul_34_17_n_7867 & mul_34_17_n_11386) | ((mul_34_17_n_7867 & mul_34_17_n_7889)
    | (mul_34_17_n_7889 & mul_34_17_n_11386)));
 assign mul_34_17_n_8611 = ((mul_34_17_n_8056 & mul_34_17_n_7439) | ((mul_34_17_n_8056 & mul_34_17_n_7669)
    | (mul_34_17_n_7669 & mul_34_17_n_7439)));
 assign mul_34_17_n_8610 = ~(mul_34_17_n_8091 ^ mul_34_17_n_7109);
 assign mul_34_17_n_8609 = ((mul_34_17_n_7893 & mul_34_17_n_8269) | ((mul_34_17_n_7893 & mul_34_17_n_7460)
    | (mul_34_17_n_7460 & mul_34_17_n_8269)));
 assign mul_34_17_n_8607 = ~(mul_34_17_n_8075 ^ mul_34_17_n_7590);
 assign mul_34_17_n_8604 = ((mul_34_17_n_7834 & mul_34_17_n_7844) | ((mul_34_17_n_7834 & mul_34_17_n_7475)
    | (mul_34_17_n_7475 & mul_34_17_n_7844)));
 assign mul_34_17_n_8602 = ((mul_34_17_n_7930 & mul_34_17_n_7845) | ((mul_34_17_n_7930 & mul_34_17_n_7984)
    | (mul_34_17_n_7984 & mul_34_17_n_7845)));
 assign mul_34_17_n_8599 = ((mul_34_17_n_7881 & mul_34_17_n_8226) | ((mul_34_17_n_7881 & mul_34_17_n_8035)
    | (mul_34_17_n_8035 & mul_34_17_n_8226)));
 assign mul_34_17_n_8598 = ~(mul_34_17_n_8100 ^ mul_34_17_n_7346);
 assign mul_34_17_n_8596 = ~(mul_34_17_n_8101 ^ mul_34_17_n_7527);
 assign mul_34_17_n_8595 = ((mul_34_17_n_206 & mul_34_17_n_11487) | ((mul_34_17_n_206 & mul_34_17_n_7666)
    | (mul_34_17_n_7666 & mul_34_17_n_11487)));
 assign mul_34_17_n_8593 = ~(mul_34_17_n_8104 ^ mul_34_17_n_7442);
 assign mul_34_17_n_8592 = ~(mul_34_17_n_8097 ^ mul_34_17_n_7448);
 assign mul_34_17_n_8550 = ~mul_34_17_n_8549;
 assign mul_34_17_n_8544 = ~mul_34_17_n_8543;
 assign mul_34_17_n_8540 = ~mul_34_17_n_8539;
 assign mul_34_17_n_8521 = ~mul_34_17_n_8520;
 assign mul_34_17_n_8518 = ~mul_34_17_n_8517;
 assign mul_34_17_n_8508 = ~mul_34_17_n_8507;
 assign mul_34_17_n_8502 = ~mul_34_17_n_8501;
 assign mul_34_17_n_8491 = ~mul_34_17_n_8492;
 assign mul_34_17_n_8490 = ~mul_34_17_n_8489;
 assign mul_34_17_n_8488 = ~mul_34_17_n_8487;
 assign mul_34_17_n_8482 = (mul_34_17_n_8002 ^ mul_34_17_n_7743);
 assign mul_34_17_n_8480 = ~(mul_34_17_n_374 | mul_34_17_n_7277);
 assign mul_34_17_n_8479 = ~(mul_34_17_n_380 | mul_34_17_n_7650);
 assign mul_34_17_n_8478 = ~(mul_34_17_n_8121 | mul_34_17_n_7645);
 assign mul_34_17_n_8477 = ~(mul_34_17_n_8134 & mul_34_17_n_7435);
 assign mul_34_17_n_8476 = ~(mul_34_17_n_8134 | mul_34_17_n_7435);
 assign mul_34_17_n_8475 = ~(mul_34_17_n_8119 | mul_34_17_n_7260);
 assign mul_34_17_n_8474 = ~(mul_34_17_n_372 | mul_34_17_n_7643);
 assign mul_34_17_n_8473 = ~(mul_34_17_n_367 | mul_34_17_n_7638);
 assign mul_34_17_n_8472 = ~(mul_34_17_n_8112 | mul_34_17_n_7657);
 assign mul_34_17_n_8574 = ~(mul_34_17_n_7887 ^ mul_34_17_n_7885);
 assign mul_34_17_n_8470 = ~(mul_34_17_n_7938 ^ mul_34_17_n_7156);
 assign mul_34_17_n_8469 = ~(mul_34_17_n_8041 ^ mul_34_17_n_166);
 assign mul_34_17_n_8468 = (mul_34_17_n_11410 ^ mul_34_17_n_11418);
 assign mul_34_17_n_8467 = ~(mul_34_17_n_378 | mul_34_17_n_7620);
 assign mul_34_17_n_8466 = ~(mul_34_17_n_8164 | mul_34_17_n_7918);
 assign mul_34_17_n_8465 = ~(mul_34_17_n_8163 | mul_34_17_n_7919);
 assign mul_34_17_n_8464 = ~(mul_34_17_n_368 | mul_34_17_n_7606);
 assign mul_34_17_n_8463 = ~(mul_34_17_n_8133 | mul_34_17_n_7424);
 assign mul_34_17_n_8462 = ~(mul_34_17_n_8133 & mul_34_17_n_7424);
 assign mul_34_17_n_8461 = ~(mul_34_17_n_8137 | mul_34_17_n_7412);
 assign mul_34_17_n_8460 = ~(mul_34_17_n_8137 & mul_34_17_n_7412);
 assign mul_34_17_n_8459 = (mul_34_17_n_11418 ^ mul_34_17_n_11410);
 assign mul_34_17_n_8458 = ~(mul_34_17_n_7843 ^ mul_34_17_n_7835);
 assign mul_34_17_n_8454 = ~(mul_34_17_n_7842 ^ mul_34_17_n_7996);
 assign mul_34_17_n_8453 = (mul_34_17_n_215 ^ mul_34_17_n_7983);
 assign mul_34_17_n_8452 = ~((mul_34_17_n_7159 | mul_34_17_n_6404) & (mul_34_17_n_8072 | mul_34_17_n_8067));
 assign mul_34_17_n_8451 = ~(mul_34_17_n_7387 ^ (mul_34_17_n_5649 ^ (mul_34_17_n_6928 ^ mul_34_17_n_5587)));
 assign mul_34_17_n_8450 = ~(mul_34_17_n_218 ^ mul_34_17_n_11470);
 assign mul_34_17_n_8449 = ~(mul_34_17_n_7895 ^ mul_34_17_n_6902);
 assign mul_34_17_n_8448 = ~((mul_34_17_n_7623 & mul_34_17_n_7436) | (mul_34_17_n_237 & mul_34_17_n_7592));
 assign mul_34_17_n_8447 = (mul_34_17_n_8044 ^ mul_34_17_n_8031);
 assign mul_34_17_n_8446 = (mul_34_17_n_11627 ^ mul_34_17_n_11631);
 assign mul_34_17_n_8445 = ~(mul_34_17_n_7941 ^ mul_34_17_n_7798);
 assign mul_34_17_n_8444 = (mul_34_17_n_8052 ^ mul_34_17_n_165);
 assign mul_34_17_n_8573 = (mul_34_17_n_7893 ^ mul_34_17_n_7460);
 assign mul_34_17_n_8443 = ~(mul_34_17_n_7913 ^ mul_34_17_n_7720);
 assign mul_34_17_n_8442 = (mul_34_17_n_11448 ^ mul_34_17_n_11392);
 assign mul_34_17_n_8441 = ~(mul_34_17_n_6940 ^ (mul_34_17_n_6247 ^ (mul_34_17_n_7157 ^ mul_34_17_n_5719)));
 assign mul_34_17_n_8572 = ~(mul_34_17_n_8015 ^ mul_34_17_n_7536);
 assign mul_34_17_n_8571 = ~(mul_34_17_n_7875 ^ mul_34_17_n_223);
 assign mul_34_17_n_8570 = ~(mul_34_17_n_11402 ^ mul_34_17_n_7685);
 assign mul_34_17_n_8440 = ~(mul_34_17_n_186 ^ mul_34_17_n_7708);
 assign mul_34_17_n_8439 = (mul_34_17_n_8022 ^ mul_34_17_n_8050);
 assign mul_34_17_n_8438 = (mul_34_17_n_7911 ^ mul_34_17_n_8016);
 assign mul_34_17_n_8437 = (mul_34_17_n_8040 ^ mul_34_17_n_8010);
 assign mul_34_17_n_8436 = ~(mul_34_17_n_8042 ^ mul_34_17_n_7707);
 assign mul_34_17_n_8435 = ~(mul_34_17_n_11382 ^ mul_34_17_n_8023);
 assign mul_34_17_n_8434 = (mul_34_17_n_11442 ^ mul_34_17_n_11440);
 assign mul_34_17_n_8433 = (mul_34_17_n_8048 ^ mul_34_17_n_7719);
 assign mul_34_17_n_8432 = ((mul_34_17_n_7739 & mul_34_17_n_7371) | ((mul_34_17_n_7739 & mul_34_17_n_7738)
    | (mul_34_17_n_7738 & mul_34_17_n_7371)));
 assign mul_34_17_n_8568 = ((mul_34_17_n_7734 & mul_34_17_n_8063) | ((mul_34_17_n_7734 & mul_34_17_n_7735)
    | (mul_34_17_n_7735 & mul_34_17_n_8063)));
 assign mul_34_17_n_8567 = ((mul_34_17_n_7714 & mul_34_17_n_11498) | ((mul_34_17_n_7714 & mul_34_17_n_185)
    | (mul_34_17_n_185 & mul_34_17_n_11498)));
 assign mul_34_17_n_8566 = ((mul_34_17_n_7459 & mul_34_17_n_7592) | ((mul_34_17_n_7459 & mul_34_17_n_7436)
    | (mul_34_17_n_7436 & mul_34_17_n_7592)));
 assign mul_34_17_n_8565 = ((mul_34_17_n_7710 & mul_34_17_n_7353) | ((mul_34_17_n_7710 & mul_34_17_n_7302)
    | (mul_34_17_n_7302 & mul_34_17_n_7353)));
 assign mul_34_17_n_8564 = ((mul_34_17_n_7501 & mul_34_17_n_7579) | ((mul_34_17_n_7501 & mul_34_17_n_7503)
    | (mul_34_17_n_7503 & mul_34_17_n_7579)));
 assign mul_34_17_n_8563 = ((mul_34_17_n_7741 & mul_34_17_n_7783) | ((mul_34_17_n_7741 & mul_34_17_n_7742)
    | (mul_34_17_n_7742 & mul_34_17_n_7783)));
 assign mul_34_17_n_8562 = ~(mul_34_17_n_8037 ^ mul_34_17_n_189);
 assign mul_34_17_n_8561 = ((mul_34_17_n_7532 & mul_34_17_n_7559) | ((mul_34_17_n_7532 & mul_34_17_n_7697)
    | (mul_34_17_n_7697 & mul_34_17_n_7559)));
 assign mul_34_17_n_8560 = ((mul_34_17_n_7599 & mul_34_17_n_7573) | ((mul_34_17_n_7599 & mul_34_17_n_7595)
    | (mul_34_17_n_7595 & mul_34_17_n_7573)));
 assign mul_34_17_n_8559 = ~(mul_34_17_n_8027 ^ mul_34_17_n_7290);
 assign mul_34_17_n_8558 = ~((mul_34_17_n_7968 & mul_34_17_n_148) | (mul_34_17_n_7976 & mul_34_17_n_6808));
 assign mul_34_17_n_8557 = ((mul_34_17_n_7740 & mul_34_17_n_7795) | ((mul_34_17_n_7740 & mul_34_17_n_7747)
    | (mul_34_17_n_7747 & mul_34_17_n_7795)));
 assign mul_34_17_n_8556 = ~(mul_34_17_n_8011 ^ mul_34_17_n_7670);
 assign mul_34_17_n_8431 = ((mul_34_17_n_7622 | mul_34_17_n_6882) & (mul_34_17_n_7971 | mul_34_17_n_7972));
 assign mul_34_17_n_8555 = ((mul_34_17_n_7670 & mul_34_17_n_7364) | ((mul_34_17_n_7670 & mul_34_17_n_7301)
    | (mul_34_17_n_7301 & mul_34_17_n_7364)));
 assign mul_34_17_n_8430 = ~(mul_34_17_n_8165 | mul_34_17_n_8070);
 assign mul_34_17_n_8554 = ((mul_34_17_n_7442 & mul_34_17_n_7379) | ((mul_34_17_n_7442 & mul_34_17_n_192)
    | (mul_34_17_n_192 & mul_34_17_n_7379)));
 assign mul_34_17_n_8553 = ~(mul_34_17_n_8001 ^ mul_34_17_n_6895);
 assign mul_34_17_n_8552 = ((mul_34_17_n_173 & mul_34_17_n_7438) | ((mul_34_17_n_173 & mul_34_17_n_7420)
    | (mul_34_17_n_7420 & mul_34_17_n_7438)));
 assign mul_34_17_n_8551 = ((mul_34_17_n_7425 & mul_34_17_n_7440) | ((mul_34_17_n_7425 & mul_34_17_n_7469)
    | (mul_34_17_n_7469 & mul_34_17_n_7440)));
 assign mul_34_17_n_8549 = ((mul_34_17_n_189 & mul_34_17_n_7375) | ((mul_34_17_n_189 & mul_34_17_n_7295)
    | (mul_34_17_n_7295 & mul_34_17_n_7375)));
 assign mul_34_17_n_8548 = ~(mul_34_17_n_8035 ^ mul_34_17_n_7881);
 assign mul_34_17_n_8547 = ((mul_34_17_n_7686 & mul_34_17_n_7351) | ((mul_34_17_n_7686 & mul_34_17_n_7695)
    | (mul_34_17_n_7695 & mul_34_17_n_7351)));
 assign mul_34_17_n_8546 = (mul_34_17_n_8069 ^ mul_34_17_n_7696);
 assign mul_34_17_n_8545 = ((mul_34_17_n_7557 & mul_34_17_n_7677) | ((mul_34_17_n_7557 & mul_34_17_n_7671)
    | (mul_34_17_n_7671 & mul_34_17_n_7677)));
 assign mul_34_17_n_8543 = ((mul_34_17_n_7730 & mul_34_17_n_7381) | ((mul_34_17_n_7730 & mul_34_17_n_7731)
    | (mul_34_17_n_7731 & mul_34_17_n_7381)));
 assign mul_34_17_n_8542 = ((mul_34_17_n_7687 & mul_34_17_n_7776) | ((mul_34_17_n_7687 & mul_34_17_n_7463)
    | (mul_34_17_n_7463 & mul_34_17_n_7776)));
 assign mul_34_17_n_8541 = ((mul_34_17_n_7500 & mul_34_17_n_7146) | ((mul_34_17_n_7500 & mul_34_17_n_6896)
    | (mul_34_17_n_6896 & mul_34_17_n_7146)));
 assign mul_34_17_n_8539 = ((mul_34_17_n_7691 & mul_34_17_n_7354) | ((mul_34_17_n_7691 & mul_34_17_n_7330)
    | (mul_34_17_n_7330 & mul_34_17_n_7354)));
 assign mul_34_17_n_8538 = ((mul_34_17_n_7544 & mul_34_17_n_7932) | ((mul_34_17_n_7544 & mul_34_17_n_7545)
    | (mul_34_17_n_7545 & mul_34_17_n_7932)));
 assign mul_34_17_n_8537 = ((mul_34_17_n_7721 & mul_34_17_n_7913) | ((mul_34_17_n_7721 & mul_34_17_n_7476)
    | (mul_34_17_n_7476 & mul_34_17_n_7913)));
 assign mul_34_17_n_8536 = ((mul_34_17_n_7467 & mul_34_17_n_7778) | ((mul_34_17_n_7467 & mul_34_17_n_7085)
    | (mul_34_17_n_7085 & mul_34_17_n_7778)));
 assign mul_34_17_n_8535 = ~(mul_34_17_n_7947 ^ mul_34_17_n_7069);
 assign mul_34_17_n_8534 = ((mul_34_17_n_7672 & mul_34_17_n_167) | ((mul_34_17_n_7672 & mul_34_17_n_162)
    | (mul_34_17_n_162 & mul_34_17_n_167)));
 assign mul_34_17_n_8533 = ((mul_34_17_n_7709 & mul_34_17_n_186) | ((mul_34_17_n_7709 & mul_34_17_n_7749)
    | (mul_34_17_n_7749 & mul_34_17_n_186)));
 assign mul_34_17_n_8532 = ((mul_34_17_n_7732 & mul_34_17_n_7767) | ((mul_34_17_n_7732 & mul_34_17_n_7733)
    | (mul_34_17_n_7733 & mul_34_17_n_7767)));
 assign mul_34_17_n_8531 = ((mul_34_17_n_7513 & mul_34_17_n_7434) | ((mul_34_17_n_7513 & mul_34_17_n_6779)
    | (mul_34_17_n_6779 & mul_34_17_n_7434)));
 assign mul_34_17_n_8530 = ((mul_34_17_n_7528 & mul_34_17_n_207) | ((mul_34_17_n_7528 & mul_34_17_n_7525)
    | (mul_34_17_n_7525 & mul_34_17_n_207)));
 assign mul_34_17_n_8529 = ((mul_34_17_n_7723 & mul_34_17_n_7363) | ((mul_34_17_n_7723 & mul_34_17_n_7725)
    | (mul_34_17_n_7725 & mul_34_17_n_7363)));
 assign mul_34_17_n_8528 = ((mul_34_17_n_7584 & mul_34_17_n_7065) | ((mul_34_17_n_7584 & mul_34_17_n_7049)
    | (mul_34_17_n_7049 & mul_34_17_n_7065)));
 assign mul_34_17_n_8527 = ((mul_34_17_n_7542 & mul_34_17_n_7058) | ((mul_34_17_n_7542 & mul_34_17_n_6454)
    | (mul_34_17_n_6454 & mul_34_17_n_7058)));
 assign mul_34_17_n_8525 = ((mul_34_17_n_7707 & mul_34_17_n_8042) | ((mul_34_17_n_7707 & mul_34_17_n_7774)
    | (mul_34_17_n_7774 & mul_34_17_n_8042)));
 assign mul_34_17_n_8524 = ~(mul_34_17_n_7953 ^ mul_34_17_n_7331);
 assign mul_34_17_n_8523 = ~(mul_34_17_n_7957 ^ mul_34_17_n_7138);
 assign mul_34_17_n_8522 = ((mul_34_17_n_7498 & mul_34_17_n_7780) | ((mul_34_17_n_7498 & mul_34_17_n_7340)
    | (mul_34_17_n_7340 & mul_34_17_n_7780)));
 assign mul_34_17_n_8520 = ((mul_34_17_n_7800 & mul_34_17_n_11500) | ((mul_34_17_n_7800 & mul_34_17_n_7799)
    | (mul_34_17_n_7799 & mul_34_17_n_11500)));
 assign mul_34_17_n_8519 = ((mul_34_17_n_7508 & mul_34_17_n_7382) | ((mul_34_17_n_7508 & mul_34_17_n_6780)
    | (mul_34_17_n_6780 & mul_34_17_n_7382)));
 assign mul_34_17_n_8517 = ((mul_34_17_n_7689 & mul_34_17_n_8046) | ((mul_34_17_n_7689 & mul_34_17_n_7690)
    | (mul_34_17_n_7690 & mul_34_17_n_8046)));
 assign mul_34_17_n_8516 = ((mul_34_17_n_7705 & mul_34_17_n_7772) | ((mul_34_17_n_7705 & mul_34_17_n_7706)
    | (mul_34_17_n_7706 & mul_34_17_n_7772)));
 assign mul_34_17_n_8515 = ((mul_34_17_n_7724 & mul_34_17_n_7779) | ((mul_34_17_n_7724 & mul_34_17_n_7511)
    | (mul_34_17_n_7511 & mul_34_17_n_7779)));
 assign mul_34_17_n_8514 = ~(mul_34_17_n_7140 ^ mul_34_17_n_7946);
 assign mul_34_17_n_8513 = ((mul_34_17_n_197 & mul_34_17_n_7566) | ((mul_34_17_n_197 & mul_34_17_n_7758)
    | (mul_34_17_n_7758 & mul_34_17_n_7566)));
 assign mul_34_17_n_8512 = ((mul_34_17_n_7696 & mul_34_17_n_7153) | ((mul_34_17_n_7696 & mul_34_17_n_7322)
    | (mul_34_17_n_7322 & mul_34_17_n_7153)));
 assign mul_34_17_n_8511 = ((mul_34_17_n_7727 & mul_34_17_n_8060) | ((mul_34_17_n_7727 & mul_34_17_n_170)
    | (mul_34_17_n_170 & mul_34_17_n_8060)));
 assign mul_34_17_n_8510 = ((mul_34_17_n_7702 & mul_34_17_n_8061) | ((mul_34_17_n_7702 & mul_34_17_n_6906)
    | (mul_34_17_n_6906 & mul_34_17_n_8061)));
 assign mul_34_17_n_8509 = ((mul_34_17_n_7587 & mul_34_17_n_7358) | ((mul_34_17_n_7587 & mul_34_17_n_7334)
    | (mul_34_17_n_7334 & mul_34_17_n_7358)));
 assign mul_34_17_n_8507 = ((mul_34_17_n_166 & mul_34_17_n_7370) | ((mul_34_17_n_166 & mul_34_17_n_6909)
    | (mul_34_17_n_6909 & mul_34_17_n_7370)));
 assign mul_34_17_n_8506 = ~(mul_34_17_n_7955 ^ mul_34_17_n_7356);
 assign mul_34_17_n_8505 = ((mul_34_17_n_7394 & mul_34_17_n_7143) | ((mul_34_17_n_7394 & mul_34_17_n_6916)
    | (mul_34_17_n_6916 & mul_34_17_n_7143)));
 assign mul_34_17_n_8504 = ((mul_34_17_n_7521 & mul_34_17_n_7149) | ((mul_34_17_n_7521 & mul_34_17_n_6911)
    | (mul_34_17_n_6911 & mul_34_17_n_7149)));
 assign mul_34_17_n_8503 = ((mul_34_17_n_191 & mul_34_17_n_7572) | ((mul_34_17_n_191 & mul_34_17_n_7424)
    | (mul_34_17_n_7424 & mul_34_17_n_7572)));
 assign mul_34_17_n_8501 = ((mul_34_17_n_7693 & mul_34_17_n_7788) | ((mul_34_17_n_7693 & mul_34_17_n_7694)
    | (mul_34_17_n_7694 & mul_34_17_n_7788)));
 assign mul_34_17_n_8500 = ((mul_34_17_n_7699 & mul_34_17_n_7771) | ((mul_34_17_n_7699 & mul_34_17_n_7317)
    | (mul_34_17_n_7317 & mul_34_17_n_7771)));
 assign mul_34_17_n_8499 = ((mul_34_17_n_7746 & mul_34_17_n_7784) | ((mul_34_17_n_7746 & mul_34_17_n_7748)
    | (mul_34_17_n_7748 & mul_34_17_n_7784)));
 assign mul_34_17_n_8498 = ((mul_34_17_n_11502 & mul_34_17_n_7346) | ((mul_34_17_n_11502 & mul_34_17_n_6913)
    | (mul_34_17_n_6913 & mul_34_17_n_7346)));
 assign mul_34_17_n_8497 = ((mul_34_17_n_7480 & mul_34_17_n_7586) | ((mul_34_17_n_7480 & mul_34_17_n_7336)
    | (mul_34_17_n_7336 & mul_34_17_n_7586)));
 assign mul_34_17_n_8496 = ~(mul_34_17_n_7956 ^ mul_34_17_n_7299);
 assign mul_34_17_n_8495 = ((mul_34_17_n_7597 & mul_34_17_n_7373) | ((mul_34_17_n_7597 & mul_34_17_n_11641)
    | (mul_34_17_n_11641 & mul_34_17_n_7373)));
 assign mul_34_17_n_8494 = ((mul_34_17_n_7796 & mul_34_17_n_11483) | ((mul_34_17_n_7796 & mul_34_17_n_7385)
    | (mul_34_17_n_7385 & mul_34_17_n_11483)));
 assign mul_34_17_n_8493 = ((mul_34_17_n_7499 & mul_34_17_n_8066) | ((mul_34_17_n_7499 & mul_34_17_n_7494)
    | (mul_34_17_n_7494 & mul_34_17_n_8066)));
 assign mul_34_17_n_8492 = ((mul_34_17_n_7763 & mul_34_17_n_7944) | ((mul_34_17_n_7763 & mul_34_17_n_156)
    | (mul_34_17_n_156 & mul_34_17_n_7944)));
 assign mul_34_17_n_8489 = ((mul_34_17_n_369 & mul_34_17_n_7552) | ((mul_34_17_n_369 & mul_34_17_n_7066)
    | (mul_34_17_n_7066 & mul_34_17_n_7552)));
 assign mul_34_17_n_8487 = ((mul_34_17_n_7711 & mul_34_17_n_7292) | ((mul_34_17_n_7711 & mul_34_17_n_6893)
    | (mul_34_17_n_6893 & mul_34_17_n_7292)));
 assign mul_34_17_n_8486 = ~(mul_34_17_n_7949 ^ mul_34_17_n_7305);
 assign mul_34_17_n_8485 = ((mul_34_17_n_7530 & mul_34_17_n_202) | ((mul_34_17_n_7530 & mul_34_17_n_7523)
    | (mul_34_17_n_7523 & mul_34_17_n_202)));
 assign mul_34_17_n_8421 = ~mul_34_17_n_247;
 assign mul_34_17_n_8414 = ~mul_34_17_n_8413;
 assign mul_34_17_n_8405 = ~mul_34_17_n_8404;
 assign mul_34_17_n_8397 = ~mul_34_17_n_8396;
 assign mul_34_17_n_8395 = ~mul_34_17_n_8394;
 assign mul_34_17_n_8391 = ~mul_34_17_n_8390;
 assign mul_34_17_n_8387 = ~mul_34_17_n_8386;
 assign mul_34_17_n_8362 = ~mul_34_17_n_8361;
 assign mul_34_17_n_8352 = ~mul_34_17_n_8353;
 assign mul_34_17_n_8335 = ~mul_34_17_n_8334;
 assign mul_34_17_n_8332 = ~mul_34_17_n_8331;
 assign mul_34_17_n_8328 = ~mul_34_17_n_8329;
 assign mul_34_17_n_8326 = ~mul_34_17_n_8327;
 assign mul_34_17_n_8324 = ~mul_34_17_n_8323;
 assign mul_34_17_n_8321 = ~(mul_34_17_n_8203 | mul_34_17_n_7608);
 assign mul_34_17_n_8314 = ((mul_34_17_n_369 | mul_34_17_n_7205) & (mul_34_17_n_242 | mul_34_17_n_7552));
 assign mul_34_17_n_8313 = ~(mul_34_17_n_7416 ^ mul_34_17_n_7855);
 assign mul_34_17_n_8312 = ~(mul_34_17_n_7984 ^ mul_34_17_n_7845);
 assign mul_34_17_n_8311 = ~(mul_34_17_n_7845 ^ mul_34_17_n_7984);
 assign mul_34_17_n_8429 = (mul_34_17_n_7887 ^ mul_34_17_n_7885);
 assign mul_34_17_n_8308 = (mul_34_17_n_7902 ^ mul_34_17_n_7751);
 assign mul_34_17_n_8307 = ~((mul_34_17_n_7768 | mul_34_17_n_6921) & (mul_34_17_n_8072 | mul_34_17_n_8068));
 assign mul_34_17_n_8305 = (mul_34_17_n_8012 ^ mul_34_17_n_11424);
 assign mul_34_17_n_8304 = (mul_34_17_n_8024 ^ mul_34_17_n_11434);
 assign mul_34_17_n_8303 = ~(mul_34_17_n_7935 ^ mul_34_17_n_158);
 assign mul_34_17_n_8302 = (mul_34_17_n_11426 ^ mul_34_17_n_8017);
 assign mul_34_17_n_8428 = ((mul_34_17_n_7598 & mul_34_17_n_7937) | ((mul_34_17_n_7598 & mul_34_17_n_6776)
    | (mul_34_17_n_6776 & mul_34_17_n_7937)));
 assign mul_34_17_n_8427 = (mul_34_17_n_11436 ^ mul_34_17_n_163);
 assign mul_34_17_n_8301 = ~((mul_34_17_n_5983 & (~mul_34_17_n_7321 & ~mul_34_17_n_6839)) | ((mul_34_17_n_5982
    & (mul_34_17_n_7321 & ~mul_34_17_n_6839)) | (mul_34_17_n_7961 & mul_34_17_n_6839)));
 assign mul_34_17_n_8300 = (mul_34_17_n_11432 ^ mul_34_17_n_11458);
 assign mul_34_17_n_8299 = (mul_34_17_n_11462 ^ mul_34_17_n_11390);
 assign mul_34_17_n_8298 = (mul_34_17_n_7538 ^ mul_34_17_n_11398);
 assign mul_34_17_n_8297 = (mul_34_17_n_229 ^ mul_34_17_n_11446);
 assign mul_34_17_n_8296 = (mul_34_17_n_8061 ^ mul_34_17_n_6906);
 assign mul_34_17_n_8426 = (mul_34_17_n_11396 ^ mul_34_17_n_11438);
 assign mul_34_17_n_8295 = (mul_34_17_n_7759 ^ mul_34_17_n_8025);
 assign mul_34_17_n_8425 = ((mul_34_17_n_7415 & mul_34_17_n_7855) | ((mul_34_17_n_7415 & mul_34_17_n_7496)
    | (mul_34_17_n_7496 & mul_34_17_n_7855)));
 assign mul_34_17_n_8294 = (mul_34_17_n_11452 ^ mul_34_17_n_11450);
 assign mul_34_17_n_8293 = (mul_34_17_n_11635 ^ mul_34_17_n_11430);
 assign mul_34_17_n_8292 = (mul_34_17_n_7880 ^ mul_34_17_n_7756);
 assign mul_34_17_n_8291 = ~(mul_34_17_n_11460 ^ mul_34_17_n_7908);
 assign mul_34_17_n_8424 = (mul_34_17_n_7867 ^ mul_34_17_n_11386);
 assign mul_34_17_n_8290 = (mul_34_17_n_7884 ^ mul_34_17_n_7903);
 assign mul_34_17_n_8423 = ((mul_34_17_n_7505 & mul_34_17_n_7919) | ((mul_34_17_n_7505 & mul_34_17_n_184)
    | (mul_34_17_n_184 & mul_34_17_n_7919)));
 assign mul_34_17_n_8289 = (mul_34_17_n_7865 ^ mul_34_17_n_11420);
 assign mul_34_17_n_8288 = (mul_34_17_n_11639 ^ mul_34_17_n_11422);
 assign mul_34_17_n_8287 = ~(mul_34_17_n_201 ^ mul_34_17_n_193);
 assign mul_34_17_n_8286 = (mul_34_17_n_11456 ^ mul_34_17_n_7926);
 assign mul_34_17_n_8285 = (mul_34_17_n_7876 ^ mul_34_17_n_7872);
 assign mul_34_17_n_8284 = (mul_34_17_n_7786 ^ mul_34_17_n_7864);
 assign mul_34_17_n_8283 = (mul_34_17_n_7882 ^ mul_34_17_n_7869);
 assign mul_34_17_n_8420 = ((mul_34_17_n_7487 & mul_34_17_n_7793) | ((mul_34_17_n_7487 & mul_34_17_n_7488)
    | (mul_34_17_n_7488 & mul_34_17_n_7793)));
 assign mul_34_17_n_8419 = ((mul_34_17_n_7489 & mul_34_17_n_7794) | ((mul_34_17_n_7489 & mul_34_17_n_7412)
    | (mul_34_17_n_7412 & mul_34_17_n_7794)));
 assign mul_34_17_n_8418 = ((mul_34_17_n_7478 & mul_34_17_n_7585) | ((mul_34_17_n_7478 & mul_34_17_n_7479)
    | (mul_34_17_n_7479 & mul_34_17_n_7585)));
 assign mul_34_17_n_8417 = ~(mul_34_17_n_7816 ^ mul_34_17_n_7090);
 assign mul_34_17_n_8416 = ((mul_34_17_n_7468 & mul_34_17_n_7588) | ((mul_34_17_n_7468 & mul_34_17_n_7423)
    | (mul_34_17_n_7423 & mul_34_17_n_7588)));
 assign mul_34_17_n_8415 = ~(mul_34_17_n_7819 ^ mul_34_17_n_7073);
 assign mul_34_17_n_8413 = ~(mul_34_17_n_7861 ^ mul_34_17_n_7430);
 assign mul_34_17_n_8412 = ((mul_34_17_n_7765 & mul_34_17_n_7590) | ((mul_34_17_n_7765 & mul_34_17_n_157)
    | (mul_34_17_n_157 & mul_34_17_n_7590)));
 assign mul_34_17_n_8411 = ((mul_34_17_n_7549 & mul_34_17_n_7555) | ((mul_34_17_n_7549 & mul_34_17_n_7311)
    | (mul_34_17_n_7311 & mul_34_17_n_7555)));
 assign mul_34_17_n_8410 = ((mul_34_17_n_193 & mul_34_17_n_8051) | ((mul_34_17_n_193 & mul_34_17_n_7312)
    | (mul_34_17_n_7312 & mul_34_17_n_8051)));
 assign mul_34_17_n_8409 = ((mul_34_17_n_7445 & mul_34_17_n_7785) | ((mul_34_17_n_7445 & mul_34_17_n_7453)
    | (mul_34_17_n_7453 & mul_34_17_n_7785)));
 assign mul_34_17_n_8408 = ~(mul_34_17_n_7820 ^ mul_34_17_n_7076);
 assign mul_34_17_n_8407 = ((mul_34_17_n_11504 & mul_34_17_n_211) | ((mul_34_17_n_11504 & mul_34_17_n_7464)
    | (mul_34_17_n_7464 & mul_34_17_n_211)));
 assign mul_34_17_n_8406 = ((mul_34_17_n_7524 & mul_34_17_n_11485) | ((mul_34_17_n_7524 & mul_34_17_n_7490)
    | (mul_34_17_n_7490 & mul_34_17_n_11485)));
 assign mul_34_17_n_8404 = ((mul_34_17_n_7539 & mul_34_17_n_7437) | ((mul_34_17_n_7539 & mul_34_17_n_6787)
    | (mul_34_17_n_6787 & mul_34_17_n_7437)));
 assign mul_34_17_n_8403 = ~((mul_34_17_n_6492 & (~mul_34_17_n_194 & ~mul_34_17_n_6915)) | ((mul_34_17_n_6491
    & (mul_34_17_n_194 & ~mul_34_17_n_6915)) | (mul_34_17_n_7963 & mul_34_17_n_6915)));
 assign mul_34_17_n_8402 = ~((mul_34_17_n_7055 & (~mul_34_17_n_7064 & ~mul_34_17_n_7506)) | ((mul_34_17_n_7054
    & (mul_34_17_n_7064 & ~mul_34_17_n_7506)) | (mul_34_17_n_7964 & mul_34_17_n_7506)));
 assign mul_34_17_n_8399 = ((mul_34_17_n_7824 & mul_34_17_n_7405) | (mul_34_17_n_7823 & mul_34_17_n_7570));
 assign mul_34_17_n_8398 = ((mul_34_17_n_7562 & mul_34_17_n_171) | ((mul_34_17_n_7562 & mul_34_17_n_199)
    | (mul_34_17_n_199 & mul_34_17_n_171)));
 assign mul_34_17_n_8396 = (mul_34_17_n_7871 ^ mul_34_17_n_7119);
 assign mul_34_17_n_8394 = ((mul_34_17_n_7533 & mul_34_17_n_7433) | ((mul_34_17_n_7533 & mul_34_17_n_7418)
    | (mul_34_17_n_7418 & mul_34_17_n_7433)));
 assign mul_34_17_n_8393 = ((mul_34_17_n_7736 & mul_34_17_n_7378) | ((mul_34_17_n_7736 & mul_34_17_n_7737)
    | (mul_34_17_n_7737 & mul_34_17_n_7378)));
 assign mul_34_17_n_8392 = ~(mul_34_17_n_7811 ^ mul_34_17_n_7145);
 assign mul_34_17_n_8390 = ((mul_34_17_n_7408 & mul_34_17_n_7679) | ((mul_34_17_n_7408 & mul_34_17_n_7534)
    | (mul_34_17_n_7534 & mul_34_17_n_7679)));
 assign mul_34_17_n_8389 = ((mul_34_17_n_7407 & mul_34_17_n_7431) | ((mul_34_17_n_7407 & mul_34_17_n_7537)
    | (mul_34_17_n_7537 & mul_34_17_n_7431)));
 assign mul_34_17_n_8388 = ((mul_34_17_n_7540 & mul_34_17_n_7556) | ((mul_34_17_n_7540 & mul_34_17_n_7550)
    | (mul_34_17_n_7550 & mul_34_17_n_7556)));
 assign mul_34_17_n_8386 = ((mul_34_17_n_7529 & mul_34_17_n_7561) | ((mul_34_17_n_7529 & mul_34_17_n_7068)
    | (mul_34_17_n_7068 & mul_34_17_n_7561)));
 assign mul_34_17_n_8385 = ((mul_34_17_n_7473 & mul_34_17_n_7057) | ((mul_34_17_n_7473 & mul_34_17_n_7050)
    | (mul_34_17_n_7050 & mul_34_17_n_7057)));
 assign mul_34_17_n_8384 = ((mul_34_17_n_7484 & mul_34_17_n_7792) | ((mul_34_17_n_7484 & mul_34_17_n_7097)
    | (mul_34_17_n_7097 & mul_34_17_n_7792)));
 assign mul_34_17_n_8383 = ((mul_34_17_n_7570 & mul_34_17_n_7060) | ((mul_34_17_n_7570 & mul_34_17_n_7053)
    | (mul_34_17_n_7053 & mul_34_17_n_7060)));
 assign mul_34_17_n_8382 = ~(mul_34_17_n_7818 ^ mul_34_17_n_7508);
 assign mul_34_17_n_8381 = ((mul_34_17_n_7455 & mul_34_17_n_11637) | ((mul_34_17_n_7455 & mul_34_17_n_7456)
    | (mul_34_17_n_7456 & mul_34_17_n_11637)));
 assign mul_34_17_n_8380 = ((mul_34_17_n_7392 & mul_34_17_n_7137) | ((mul_34_17_n_7392 & mul_34_17_n_7391)
    | (mul_34_17_n_7391 & mul_34_17_n_7137)));
 assign mul_34_17_n_8379 = ((mul_34_17_n_7491 & mul_34_17_n_7056) | ((mul_34_17_n_7491 & mul_34_17_n_7051)
    | (mul_34_17_n_7051 & mul_34_17_n_7056)));
 assign mul_34_17_n_8378 = ((mul_34_17_n_7531 & mul_34_17_n_7766) | ((mul_34_17_n_7531 & mul_34_17_n_7313)
    | (mul_34_17_n_7313 & mul_34_17_n_7766)));
 assign mul_34_17_n_8377 = ~(mul_34_17_n_7808 ^ mul_34_17_n_7376);
 assign mul_34_17_n_8376 = ((mul_34_17_n_7546 & mul_34_17_n_7128) | ((mul_34_17_n_7546 & mul_34_17_n_7547)
    | (mul_34_17_n_7547 & mul_34_17_n_7128)));
 assign mul_34_17_n_8375 = ((mul_34_17_n_7548 & mul_34_17_n_7782) | ((mul_34_17_n_7548 & mul_34_17_n_7109)
    | (mul_34_17_n_7109 & mul_34_17_n_7782)));
 assign mul_34_17_n_8374 = ((mul_34_17_n_7450 & mul_34_17_n_7129) | ((mul_34_17_n_7450 & mul_34_17_n_7451)
    | (mul_34_17_n_7451 & mul_34_17_n_7129)));
 assign mul_34_17_n_8373 = ((mul_34_17_n_7461 & mul_34_17_n_7791) | ((mul_34_17_n_7461 & mul_34_17_n_7507)
    | (mul_34_17_n_7507 & mul_34_17_n_7791)));
 assign mul_34_17_n_8372 = ~(mul_34_17_n_7958 ^ mul_34_17_n_7121);
 assign mul_34_17_n_8371 = ((mul_34_17_n_7465 & mul_34_17_n_7591) | ((mul_34_17_n_7465 & mul_34_17_n_7466)
    | (mul_34_17_n_7466 & mul_34_17_n_7591)));
 assign mul_34_17_n_8370 = ((mul_34_17_n_7514 & mul_34_17_n_168) | ((mul_34_17_n_7514 & mul_34_17_n_7516)
    | (mul_34_17_n_7516 & mul_34_17_n_168)));
 assign mul_34_17_n_8369 = ((mul_34_17_n_161 & mul_34_17_n_7553) | ((mul_34_17_n_161 & mul_34_17_n_7309)
    | (mul_34_17_n_7309 & mul_34_17_n_7553)));
 assign mul_34_17_n_8368 = ((mul_34_17_n_7393 & mul_34_17_n_7806) | ((mul_34_17_n_7393 & mul_34_17_n_7427)
    | (mul_34_17_n_7427 & mul_34_17_n_7806)));
 assign mul_34_17_n_8282 = ~(mul_34_17_n_7939 ^ mul_34_17_n_7383);
 assign mul_34_17_n_8367 = ~(mul_34_17_n_7158 ^ (mul_34_17_n_5530 ^ (mul_34_17_n_6805 ^ mul_34_17_n_5538)));
 assign mul_34_17_n_8366 = ((mul_34_17_n_7495 & mul_34_17_n_7580) | ((mul_34_17_n_7495 & mul_34_17_n_7704)
    | (mul_34_17_n_7704 & mul_34_17_n_7580)));
 assign mul_34_17_n_8365 = ((mul_34_17_n_7413 & mul_34_17_n_7682) | ((mul_34_17_n_7413 & mul_34_17_n_7517)
    | (mul_34_17_n_7517 & mul_34_17_n_7682)));
 assign mul_34_17_n_8364 = ((mul_34_17_n_7675 & mul_34_17_n_7441) | ((mul_34_17_n_7675 & mul_34_17_n_7493)
    | (mul_34_17_n_7493 & mul_34_17_n_7441)));
 assign mul_34_17_n_8363 = ((mul_34_17_n_7472 & mul_34_17_n_7935) | ((mul_34_17_n_7472 & mul_34_17_n_7470)
    | (mul_34_17_n_7470 & mul_34_17_n_7935)));
 assign mul_34_17_n_8361 = ((mul_34_17_n_7698 & mul_34_17_n_11633) | ((mul_34_17_n_7698 & mul_34_17_n_7760)
    | (mul_34_17_n_7760 & mul_34_17_n_11633)));
 assign mul_34_17_n_8360 = ((mul_34_17_n_7509 & mul_34_17_n_11492) | ((mul_34_17_n_7509 & mul_34_17_n_7316)
    | (mul_34_17_n_7316 & mul_34_17_n_11492)));
 assign mul_34_17_n_8359 = ((mul_34_17_n_169 & mul_34_17_n_7123) | ((mul_34_17_n_169 & mul_34_17_n_7447)
    | (mul_34_17_n_7447 & mul_34_17_n_7123)));
 assign mul_34_17_n_8358 = ((mul_34_17_n_7506 & mul_34_17_n_7064) | ((mul_34_17_n_7506 & mul_34_17_n_7054)
    | (mul_34_17_n_7054 & mul_34_17_n_7064)));
 assign mul_34_17_n_8357 = ~(mul_34_17_n_7821 ^ mul_34_17_n_7368);
 assign mul_34_17_n_8356 = ((mul_34_17_n_7769 & mul_34_17_n_7678) | ((mul_34_17_n_7769 & mul_34_17_n_6894)
    | (mul_34_17_n_6894 & mul_34_17_n_7678)));
 assign mul_34_17_n_8355 = ~(mul_34_17_n_7813 ^ mul_34_17_n_178);
 assign mul_34_17_n_8354 = ~(mul_34_17_n_7337 ^ mul_34_17_n_7814);
 assign mul_34_17_n_8353 = (mul_34_17_n_7936 ^ mul_34_17_n_7350);
 assign mul_34_17_n_8349 = ~(mul_34_17_n_7810 ^ mul_34_17_n_7113);
 assign mul_34_17_n_8348 = ((mul_34_17_n_5510 & (~mul_34_17_n_6907 & ~mul_34_17_n_7954)) | ((mul_34_17_n_5511
    & (mul_34_17_n_6907 & ~mul_34_17_n_7954)) | (mul_34_17_n_7587 & mul_34_17_n_7954)));
 assign mul_34_17_n_8346 = ((mul_34_17_n_7395 & mul_34_17_n_7577) | ((mul_34_17_n_7395 & mul_34_17_n_7396)
    | (mul_34_17_n_7396 & mul_34_17_n_7577)));
 assign mul_34_17_n_8344 = ((mul_34_17_n_7486 & mul_34_17_n_7581) | ((mul_34_17_n_7486 & mul_34_17_n_7091)
    | (mul_34_17_n_7091 & mul_34_17_n_7581)));
 assign mul_34_17_n_8343 = ~((mul_34_17_n_5876 & (~mul_34_17_n_6796 & ~mul_34_17_n_7812)) | ((mul_34_17_n_5875
    & (mul_34_17_n_6796 & ~mul_34_17_n_7812)) | (mul_34_17_n_7563 & mul_34_17_n_7812)));
 assign mul_34_17_n_8342 = ~(mul_34_17_n_7815 ^ mul_34_17_n_7070);
 assign mul_34_17_n_8341 = ((mul_34_17_n_7446 & mul_34_17_n_7560) | ((mul_34_17_n_7446 & mul_34_17_n_7449)
    | (mul_34_17_n_7449 & mul_34_17_n_7560)));
 assign mul_34_17_n_8281 = (mul_34_17_n_7942 ^ mul_34_17_n_7787);
 assign mul_34_17_n_8340 = ((mul_34_17_n_7715 & mul_34_17_n_7775) | ((mul_34_17_n_7715 & mul_34_17_n_7718)
    | (mul_34_17_n_7718 & mul_34_17_n_7775)));
 assign mul_34_17_n_8339 = ((mul_34_17_n_7482 & mul_34_17_n_7582) | ((mul_34_17_n_7482 & mul_34_17_n_7087)
    | (mul_34_17_n_7087 & mul_34_17_n_7582)));
 assign mul_34_17_n_8338 = ((mul_34_17_n_7444 & mul_34_17_n_7568) | ((mul_34_17_n_7444 & mul_34_17_n_7443)
    | (mul_34_17_n_7443 & mul_34_17_n_7568)));
 assign mul_34_17_n_8337 = ((mul_34_17_n_7713 & mul_34_17_n_7770) | ((mul_34_17_n_7713 & mul_34_17_n_7458)
    | (mul_34_17_n_7458 & mul_34_17_n_7770)));
 assign mul_34_17_n_8336 = ((mul_34_17_n_7527 & mul_34_17_n_7564) | ((mul_34_17_n_7527 & mul_34_17_n_7526)
    | (mul_34_17_n_7526 & mul_34_17_n_7564)));
 assign mul_34_17_n_8334 = ((mul_34_17_n_7522 & mul_34_17_n_7567) | ((mul_34_17_n_7522 & mul_34_17_n_181)
    | (mul_34_17_n_181 & mul_34_17_n_7567)));
 assign mul_34_17_n_8333 = ((mul_34_17_n_7512 & mul_34_17_n_7905) | ((mul_34_17_n_7512 & mul_34_17_n_7688)
    | (mul_34_17_n_7688 & mul_34_17_n_7905)));
 assign mul_34_17_n_8331 = ~(mul_34_17_n_7143 ^ (mul_34_17_n_6916 ^ (mul_34_17_n_6803 ^ mul_34_17_n_5552)));
 assign mul_34_17_n_8330 = ((mul_34_17_n_7722 & mul_34_17_n_11496) | ((mul_34_17_n_7722 & mul_34_17_n_7518)
    | (mul_34_17_n_7518 & mul_34_17_n_11496)));
 assign mul_34_17_n_8329 = ~(mul_34_17_n_7948 ^ mul_34_17_n_7082);
 assign mul_34_17_n_8327 = ~(mul_34_17_n_7521 ^ mul_34_17_n_7950);
 assign mul_34_17_n_8325 = ((mul_34_17_n_7481 & mul_34_17_n_7777) | ((mul_34_17_n_7481 & mul_34_17_n_7726)
    | (mul_34_17_n_7726 & mul_34_17_n_7777)));
 assign mul_34_17_n_8323 = ~(mul_34_17_n_7940 ^ mul_34_17_n_7103);
 assign mul_34_17_n_8271 = ~mul_34_17_n_8270;
 assign mul_34_17_n_8258 = ~mul_34_17_n_8257;
 assign mul_34_17_n_8249 = ~mul_34_17_n_8250;
 assign mul_34_17_n_8244 = ~mul_34_17_n_8243;
 assign mul_34_17_n_8239 = ~mul_34_17_n_8238;
 assign mul_34_17_n_8230 = ~mul_34_17_n_8229;
 assign mul_34_17_n_8222 = ~(mul_34_17_n_8072 | mul_34_17_n_8067);
 assign mul_34_17_n_8221 = ~(mul_34_17_n_375 | mul_34_17_n_6450);
 assign mul_34_17_n_8220 = ~(mul_34_17_n_8037 & mul_34_17_n_189);
 assign mul_34_17_n_8219 = ~(mul_34_17_n_8037 | mul_34_17_n_189);
 assign mul_34_17_n_8218 = (mul_34_17_n_7689 ^ mul_34_17_n_7690);
 assign mul_34_17_n_8217 = ~(mul_34_17_n_221 & mul_34_17_n_7754);
 assign mul_34_17_n_8216 = ~(mul_34_17_n_7842 & mul_34_17_n_7996);
 assign mul_34_17_n_8215 = ~(mul_34_17_n_8026 | mul_34_17_n_7290);
 assign mul_34_17_n_8214 = ~(mul_34_17_n_8027 | mul_34_17_n_7289);
 assign mul_34_17_n_8213 = ~(mul_34_17_n_8001 & mul_34_17_n_6895);
 assign mul_34_17_n_8212 = ~(mul_34_17_n_8001 | mul_34_17_n_6895);
 assign mul_34_17_n_8210 = ~(mul_34_17_n_213 | mul_34_17_n_7978);
 assign mul_34_17_n_8209 = ~(mul_34_17_n_7528 ^ mul_34_17_n_7525);
 assign mul_34_17_n_8280 = ~(mul_34_17_n_7901 & mul_34_17_n_7750);
 assign mul_34_17_n_8208 = ~(mul_34_17_n_7768 | (mul_34_17_n_6815 | (mul_34_17_n_7803 | mul_34_17_n_7366)));
 assign mul_34_17_n_8207 = ~(mul_34_17_n_7937 | mul_34_17_n_249);
 assign mul_34_17_n_8206 = ~(mul_34_17_n_8011 & mul_34_17_n_7670);
 assign mul_34_17_n_8205 = ~(mul_34_17_n_8011 | mul_34_17_n_7670);
 assign mul_34_17_n_8204 = ~(mul_34_17_n_377 | mul_34_17_n_7247);
 assign mul_34_17_n_8203 = (mul_34_17_n_7763 ^ mul_34_17_n_156);
 assign mul_34_17_n_8202 = ~((mul_34_17_n_7216 & mul_34_17_n_6476) | (mul_34_17_n_7661 & mul_34_17_n_7294));
 assign mul_34_17_n_8201 = ~(mul_34_17_n_7673 ^ mul_34_17_n_167);
 assign mul_34_17_n_8200 = ((mul_34_17_n_6910 | mul_34_17_n_5514) & (mul_34_17_n_7703 | mul_34_17_n_155));
 assign mul_34_17_n_8199 = ~(mul_34_17_n_6930 ^ (mul_34_17_n_6028 ^ (mul_34_17_n_6929 ^ mul_34_17_n_6031)));
 assign mul_34_17_n_8197 = ~(mul_34_17_n_7796 ^ mul_34_17_n_7385);
 assign mul_34_17_n_8279 = ~(mul_34_17_n_8067 & mul_34_17_n_8068);
 assign mul_34_17_n_8196 = ~(mul_34_17_n_7800 ^ mul_34_17_n_7799);
 assign mul_34_17_n_8195 = ~(mul_34_17_n_7594 ^ mul_34_17_n_7797);
 assign mul_34_17_n_8278 = (mul_34_17_n_7758 ^ mul_34_17_n_197);
 assign mul_34_17_n_8194 = (mul_34_17_n_7686 ^ mul_34_17_n_7351);
 assign mul_34_17_n_8193 = (mul_34_17_n_7597 ^ mul_34_17_n_11641);
 assign mul_34_17_n_8192 = (mul_34_17_n_7747 ^ mul_34_17_n_7740);
 assign mul_34_17_n_8277 = ~((mul_34_17_n_382 & mul_34_17_n_6645) | (mul_34_17_n_7655 & mul_34_17_n_5853));
 assign mul_34_17_n_8191 = (mul_34_17_n_7699 ^ mul_34_17_n_7771);
 assign mul_34_17_n_8190 = (mul_34_17_n_7698 ^ mul_34_17_n_7760);
 assign mul_34_17_n_8189 = (mul_34_17_n_7559 ^ mul_34_17_n_7532);
 assign mul_34_17_n_8188 = ~(mul_34_17_n_7901 | mul_34_17_n_7750);
 assign mul_34_17_n_8187 = ~(mul_34_17_n_7631 & (mul_34_17_n_7632 & (mul_34_17_n_7804 & mul_34_17_n_6935)));
 assign mul_34_17_n_8186 = ~(mul_34_17_n_6932 ^ (mul_34_17_n_6033 ^ (mul_34_17_n_6925 ^ mul_34_17_n_6071)));
 assign mul_34_17_n_8185 = ~(mul_34_17_n_7599 ^ mul_34_17_n_7595);
 assign mul_34_17_n_8184 = (mul_34_17_n_7354 ^ mul_34_17_n_7691);
 assign mul_34_17_n_8276 = (mul_34_17_n_7693 ^ mul_34_17_n_7694);
 assign mul_34_17_n_8183 = (mul_34_17_n_7741 ^ mul_34_17_n_7742);
 assign mul_34_17_n_8182 = (mul_34_17_n_7715 ^ mul_34_17_n_7775);
 assign mul_34_17_n_8181 = (mul_34_17_n_7529 ^ mul_34_17_n_7561);
 assign mul_34_17_n_8275 = (mul_34_17_n_7732 ^ mul_34_17_n_7733);
 assign mul_34_17_n_8180 = (mul_34_17_n_169 ^ mul_34_17_n_7447);
 assign mul_34_17_n_8179 = (mul_34_17_n_7784 ^ mul_34_17_n_7746);
 assign mul_34_17_n_8178 = ~(mul_34_17_n_11490 ^ mul_34_17_n_7603);
 assign mul_34_17_n_8177 = ~(mul_34_17_n_7887 & mul_34_17_n_7885);
 assign mul_34_17_n_8176 = (mul_34_17_n_7723 ^ mul_34_17_n_7725);
 assign mul_34_17_n_8175 = (mul_34_17_n_7381 ^ mul_34_17_n_7730);
 assign mul_34_17_n_8274 = ((mul_34_17_n_6781 & mul_34_17_n_7589) | ((mul_34_17_n_6781 & mul_34_17_n_27)
    | (mul_34_17_n_27 & mul_34_17_n_7589)));
 assign mul_34_17_n_8174 = (mul_34_17_n_7445 ^ mul_34_17_n_7785);
 assign mul_34_17_n_8273 = (mul_34_17_n_7738 ^ mul_34_17_n_7371);
 assign mul_34_17_n_8272 = ~(mul_34_17_n_7625 & (mul_34_17_n_7627 & (mul_34_17_n_6872 & mul_34_17_n_6438)));
 assign mul_34_17_n_8270 = ((mul_34_17_n_178 & mul_34_17_n_7127) | ((mul_34_17_n_178 & mul_34_17_n_59)
    | (mul_34_17_n_59 & mul_34_17_n_7127)));
 assign mul_34_17_n_8269 = ((mul_34_17_n_7300 & mul_34_17_n_7362) | ((mul_34_17_n_7300 & mul_34_17_n_176)
    | (mul_34_17_n_176 & mul_34_17_n_7362)));
 assign mul_34_17_n_8268 = ~(mul_34_17_n_7401 ^ mul_34_17_n_7297);
 assign mul_34_17_n_8267 = ((mul_34_17_n_7335 & mul_34_17_n_7355) | ((mul_34_17_n_7335 & mul_34_17_n_7332)
    | (mul_34_17_n_7332 & mul_34_17_n_7355)));
 assign mul_34_17_n_8266 = ((mul_34_17_n_7280 & mul_34_17_n_150) | (mul_34_17_n_7630 & mul_34_17_n_6448));
 assign mul_34_17_n_8265 = ((mul_34_17_n_7076 & mul_34_17_n_6802) | ((mul_34_17_n_7076 & mul_34_17_n_7304)
    | (mul_34_17_n_7304 & mul_34_17_n_6802)));
 assign mul_34_17_n_8264 = ~((mul_34_17_n_381 & mul_34_17_n_6643) | (mul_34_17_n_7656 & mul_34_17_n_5855));
 assign mul_34_17_n_8263 = ((mul_34_17_n_7250 & mul_34_17_n_6924) | (mul_34_17_n_7618 & mul_34_17_n_6435));
 assign mul_34_17_n_8262 = ((mul_34_17_n_7327 & mul_34_17_n_7349) | ((mul_34_17_n_7327 & mul_34_17_n_11643)
    | (mul_34_17_n_11643 & mul_34_17_n_7349)));
 assign mul_34_17_n_8261 = ((mul_34_17_n_7324 & mul_34_17_n_7357) | ((mul_34_17_n_7324 & mul_34_17_n_7323)
    | (mul_34_17_n_7323 & mul_34_17_n_7357)));
 assign mul_34_17_n_8260 = ((mul_34_17_n_7219 & mul_34_17_n_7238) | (mul_34_17_n_7660 & mul_34_17_n_7165));
 assign mul_34_17_n_8259 = ((mul_34_17_n_7090 & mul_34_17_n_7135) | ((mul_34_17_n_7090 & mul_34_17_n_5707)
    | (mul_34_17_n_5707 & mul_34_17_n_7135)));
 assign mul_34_17_n_8257 = ((mul_34_17_n_7333 & mul_34_17_n_7367) | ((mul_34_17_n_7333 & mul_34_17_n_7337)
    | (mul_34_17_n_7337 & mul_34_17_n_7367)));
 assign mul_34_17_n_8256 = ((mul_34_17_n_7209 & mul_34_17_n_6662) | (mul_34_17_n_7662 & mul_34_17_n_5836));
 assign mul_34_17_n_8255 = ((mul_34_17_n_7338 & mul_34_17_n_7145) | ((mul_34_17_n_7338 & mul_34_17_n_11520)
    | (mul_34_17_n_11520 & mul_34_17_n_7145)));
 assign mul_34_17_n_8254 = ((mul_34_17_n_7092 & mul_34_17_n_7430) | ((mul_34_17_n_7092 & mul_34_17_n_7072)
    | (mul_34_17_n_7072 & mul_34_17_n_7430)));
 assign mul_34_17_n_8253 = ((mul_34_17_n_7293 & mul_34_17_n_7305) | ((mul_34_17_n_7293 & mul_34_17_n_6477)
    | (mul_34_17_n_6477 & mul_34_17_n_7305)));
 assign mul_34_17_n_8252 = ~(mul_34_17_n_7605 ^ mul_34_17_n_7360);
 assign mul_34_17_n_8250 = ~((mul_34_17_n_388 & mul_34_17_n_6409) | (mul_34_17_n_7619 & mul_34_17_n_5868));
 assign mul_34_17_n_8248 = ((mul_34_17_n_385 & mul_34_17_n_6807) | (mul_34_17_n_7629 & mul_34_17_n_6439));
 assign mul_34_17_n_8247 = ((mul_34_17_n_6603 & mul_34_17_n_7565) | ((mul_34_17_n_6603 & mul_34_17_n_6908)
    | (mul_34_17_n_6908 & mul_34_17_n_7565)));
 assign mul_34_17_n_8246 = ((mul_34_17_n_7106 & mul_34_17_n_386) | ((mul_34_17_n_7106 & mul_34_17_n_7095)
    | (mul_34_17_n_7095 & mul_34_17_n_386)));
 assign mul_34_17_n_8245 = ~(mul_34_17_n_7600 ^ mul_34_17_n_7345);
 assign mul_34_17_n_8243 = ((mul_34_17_n_7105 & mul_34_17_n_7787) | ((mul_34_17_n_7105 & mul_34_17_n_6331)
    | (mul_34_17_n_6331 & mul_34_17_n_7787)));
 assign mul_34_17_n_8242 = ((mul_34_17_n_7099 & mul_34_17_n_7125) | ((mul_34_17_n_7099 & mul_34_17_n_7070)
    | (mul_34_17_n_7070 & mul_34_17_n_7125)));
 assign mul_34_17_n_8241 = ((mul_34_17_n_379 & mul_34_17_n_6685) | (mul_34_17_n_7642 & mul_34_17_n_6122));
 assign mul_34_17_n_8240 = ((mul_34_17_n_7100 & mul_34_17_n_7593) | ((mul_34_17_n_7100 & mul_34_17_n_7118)
    | (mul_34_17_n_7118 & mul_34_17_n_7593)));
 assign mul_34_17_n_8238 = ((mul_34_17_n_7331 & mul_34_17_n_7359) | ((mul_34_17_n_7331 & mul_34_17_n_6778)
    | (mul_34_17_n_6778 & mul_34_17_n_7359)));
 assign mul_34_17_n_8237 = ((mul_34_17_n_7115 & mul_34_17_n_183) | ((mul_34_17_n_7115 & mul_34_17_n_7116)
    | (mul_34_17_n_7116 & mul_34_17_n_183)));
 assign mul_34_17_n_8236 = ((mul_34_17_n_7289 & mul_34_17_n_7348) | ((mul_34_17_n_7289 & mul_34_17_n_5944)
    | (mul_34_17_n_5944 & mul_34_17_n_7348)));
 assign mul_34_17_n_8235 = ((mul_34_17_n_7191 & mul_34_17_n_6652) | (mul_34_17_n_7628 & mul_34_17_n_5867));
 assign mul_34_17_n_8234 = ((mul_34_17_n_7069 & mul_34_17_n_7377) | ((mul_34_17_n_7069 & mul_34_17_n_6901)
    | (mul_34_17_n_6901 & mul_34_17_n_7377)));
 assign mul_34_17_n_8233 = ~(mul_34_17_n_7604 ^ mul_34_17_n_7344);
 assign mul_34_17_n_8232 = ((mul_34_17_n_7339 & mul_34_17_n_7554) | ((mul_34_17_n_7339 & mul_34_17_n_7071)
    | (mul_34_17_n_7071 & mul_34_17_n_7554)));
 assign mul_34_17_n_8231 = ((mul_34_17_n_198 & mul_34_17_n_7380) | ((mul_34_17_n_198 & mul_34_17_n_7307)
    | (mul_34_17_n_7307 & mul_34_17_n_7380)));
 assign mul_34_17_n_8229 = ((mul_34_17_n_7113 & mul_34_17_n_7120) | ((mul_34_17_n_7113 & mul_34_17_n_7077)
    | (mul_34_17_n_7077 & mul_34_17_n_7120)));
 assign mul_34_17_n_8228 = ((mul_34_17_n_383 & mul_34_17_n_6684) | (mul_34_17_n_7665 & mul_34_17_n_5863));
 assign mul_34_17_n_8227 = ((mul_34_17_n_7329 & mul_34_17_n_7140) | ((mul_34_17_n_7329 & mul_34_17_n_6575)
    | (mul_34_17_n_6575 & mul_34_17_n_7140)));
 assign mul_34_17_n_8226 = ((mul_34_17_n_7079 & mul_34_17_n_6808) | ((mul_34_17_n_7079 & mul_34_17_n_7310)
    | (mul_34_17_n_7310 & mul_34_17_n_6808)));
 assign mul_34_17_n_8224 = ((mul_34_17_n_7075 & mul_34_17_n_6798) | ((mul_34_17_n_7075 & mul_34_17_n_6340)
    | (mul_34_17_n_6340 & mul_34_17_n_6798)));
 assign mul_34_17_n_8223 = ((mul_34_17_n_7267 & mul_34_17_n_6926) | (mul_34_17_n_7652 & mul_34_17_n_6444));
 assign mul_34_17_n_8164 = ~mul_34_17_n_8163;
 assign mul_34_17_n_8155 = ~mul_34_17_n_8154;
 assign mul_34_17_n_8147 = ~mul_34_17_n_8146;
 assign mul_34_17_n_8128 = ~mul_34_17_n_8127;
 assign mul_34_17_n_8123 = ~(mul_34_17_n_7414 ^ mul_34_17_n_7684);
 assign mul_34_17_n_8121 = ~(mul_34_17_n_6810 ^ (mul_34_17_n_5582 ^ (mul_34_17_n_6811 ^ mul_34_17_n_5574)));
 assign mul_34_17_n_8120 = (mul_34_17_n_7677 ^ mul_34_17_n_7671);
 assign mul_34_17_n_8119 = (mul_34_17_n_7671 ^ mul_34_17_n_7677);
 assign mul_34_17_n_8118 = ~(mul_34_17_n_373 | mul_34_17_n_7263);
 assign mul_34_17_n_8115 = (mul_34_17_n_156 ^ mul_34_17_n_7763);
 assign mul_34_17_n_8113 = ~(mul_34_17_n_11487 ^ mul_34_17_n_7666);
 assign mul_34_17_n_8112 = ~(mul_34_17_n_7666 ^ mul_34_17_n_11487);
 assign mul_34_17_n_8108 = ~(mul_34_17_n_7441 ^ mul_34_17_n_7675);
 assign mul_34_17_n_8173 = (mul_34_17_n_7778 ^ mul_34_17_n_7467);
 assign mul_34_17_n_8106 = (mul_34_17_n_7550 ^ mul_34_17_n_7540);
 assign mul_34_17_n_8105 = (mul_34_17_n_7706 ^ mul_34_17_n_7772);
 assign mul_34_17_n_8104 = (mul_34_17_n_192 ^ mul_34_17_n_7379);
 assign mul_34_17_n_8172 = (mul_34_17_n_7530 ^ mul_34_17_n_7523);
 assign mul_34_17_n_8171 = (mul_34_17_n_369 ^ mul_34_17_n_7552);
 assign mul_34_17_n_8103 = ~(mul_34_17_n_7586 ^ mul_34_17_n_7480);
 assign mul_34_17_n_8102 = (mul_34_17_n_7687 ^ mul_34_17_n_7776);
 assign mul_34_17_n_8101 = (mul_34_17_n_7564 ^ mul_34_17_n_7526);
 assign mul_34_17_n_8100 = (mul_34_17_n_11502 ^ mul_34_17_n_6913);
 assign mul_34_17_n_8099 = (mul_34_17_n_7450 ^ mul_34_17_n_7451);
 assign mul_34_17_n_8098 = (mul_34_17_n_11485 ^ mul_34_17_n_7524);
 assign mul_34_17_n_8097 = (mul_34_17_n_7560 ^ mul_34_17_n_7446);
 assign mul_34_17_n_8096 = (mul_34_17_n_11492 ^ mul_34_17_n_7509);
 assign mul_34_17_n_8095 = ~(mul_34_17_n_6806 ^ (mul_34_17_n_5586 ^ (mul_34_17_n_6809 ^ mul_34_17_n_5620)));
 assign mul_34_17_n_8094 = (mul_34_17_n_7553 ^ mul_34_17_n_161);
 assign mul_34_17_n_8093 = (mul_34_17_n_7737 ^ mul_34_17_n_7736);
 assign mul_34_17_n_8092 = (mul_34_17_n_7531 ^ mul_34_17_n_7313);
 assign mul_34_17_n_8091 = (mul_34_17_n_7548 ^ mul_34_17_n_7782);
 assign mul_34_17_n_8090 = (mul_34_17_n_7710 ^ mul_34_17_n_7353);
 assign mul_34_17_n_8170 = (mul_34_17_n_11496 ^ mul_34_17_n_7722);
 assign mul_34_17_n_8089 = (mul_34_17_n_7458 ^ mul_34_17_n_7770);
 assign mul_34_17_n_8088 = (mul_34_17_n_7688 ^ mul_34_17_n_7512);
 assign mul_34_17_n_8169 = (mul_34_17_n_168 ^ mul_34_17_n_7516);
 assign mul_34_17_n_8087 = (mul_34_17_n_7461 ^ mul_34_17_n_7507);
 assign mul_34_17_n_8168 = (mul_34_17_n_7522 ^ mul_34_17_n_181);
 assign mul_34_17_n_8167 = (mul_34_17_n_7455 ^ mul_34_17_n_7456);
 assign mul_34_17_n_8086 = (mul_34_17_n_7714 ^ mul_34_17_n_185);
 assign mul_34_17_n_8166 = ~(mul_34_17_n_170 ^ mul_34_17_n_7727);
 assign mul_34_17_n_8165 = ~(mul_34_17_n_7589 ^ mul_34_17_n_7596);
 assign mul_34_17_n_8085 = (mul_34_17_n_7546 ^ mul_34_17_n_7547);
 assign mul_34_17_n_8084 = (mul_34_17_n_7443 ^ mul_34_17_n_7444);
 assign mul_34_17_n_8163 = ~(mul_34_17_n_7504 ^ mul_34_17_n_184);
 assign mul_34_17_n_8162 = (mul_34_17_n_7498 ^ mul_34_17_n_7340);
 assign mul_34_17_n_8083 = (mul_34_17_n_7580 ^ mul_34_17_n_7495);
 assign mul_34_17_n_8082 = (mul_34_17_n_7549 ^ mul_34_17_n_7311);
 assign mul_34_17_n_8161 = (mul_34_17_n_5514 ^ mul_34_17_n_7703);
 assign mul_34_17_n_8160 = (mul_34_17_n_6910 ^ mul_34_17_n_155);
 assign mul_34_17_n_8081 = (mul_34_17_n_7554 ^ mul_34_17_n_7071);
 assign mul_34_17_n_8080 = (mul_34_17_n_7484 ^ mul_34_17_n_7792);
 assign mul_34_17_n_8079 = (mul_34_17_n_7488 ^ mul_34_17_n_7487);
 assign mul_34_17_n_8078 = (mul_34_17_n_7581 ^ mul_34_17_n_7486);
 assign mul_34_17_n_8077 = (mul_34_17_n_7582 ^ mul_34_17_n_7482);
 assign mul_34_17_n_8076 = (mul_34_17_n_7466 ^ mul_34_17_n_7591);
 assign mul_34_17_n_8159 = (mul_34_17_n_7459 ^ mul_34_17_n_7436);
 assign mul_34_17_n_8075 = (mul_34_17_n_157 ^ mul_34_17_n_7765);
 assign mul_34_17_n_8074 = (mul_34_17_n_7478 ^ mul_34_17_n_7479);
 assign mul_34_17_n_8073 = (mul_34_17_n_7777 ^ mul_34_17_n_7481);
 assign mul_34_17_n_8158 = ((mul_34_17_n_6794 & mul_34_17_n_7122) | ((mul_34_17_n_6794 & mul_34_17_n_7078)
    | (mul_34_17_n_7078 & mul_34_17_n_7122)));
 assign mul_34_17_n_8157 = ((mul_34_17_n_7308 & mul_34_17_n_7376) | ((mul_34_17_n_7308 & mul_34_17_n_6616)
    | (mul_34_17_n_6616 & mul_34_17_n_7376)));
 assign mul_34_17_n_8156 = ((mul_34_17_n_7320 & mul_34_17_n_6649) | ((mul_34_17_n_7320 & mul_34_17_n_6895)
    | (mul_34_17_n_6895 & mul_34_17_n_6649)));
 assign mul_34_17_n_8154 = ~((mul_34_17_n_6967 & mul_34_17_n_6362) | (mul_34_17_n_7644 & mul_34_17_n_6123));
 assign mul_34_17_n_8153 = ~(mul_34_17_n_7397 ^ mul_34_17_n_7155);
 assign mul_34_17_n_8152 = ((mul_34_17_n_7028 & mul_34_17_n_6390) | (mul_34_17_n_7647 & mul_34_17_n_5832));
 assign mul_34_17_n_8151 = ((mul_34_17_n_187 & mul_34_17_n_7369) | ((mul_34_17_n_187 & mul_34_17_n_6914)
    | (mul_34_17_n_6914 & mul_34_17_n_7369)));
 assign mul_34_17_n_8150 = ~((mul_34_17_n_6604 & (~mul_34_17_n_6908 & ~mul_34_17_n_7565)) | ((mul_34_17_n_6603
    & (mul_34_17_n_6908 & ~mul_34_17_n_7565)) | (mul_34_17_n_7403 & mul_34_17_n_7565)));
 assign mul_34_17_n_8149 = ((mul_34_17_n_7101 & mul_34_17_n_7154) | ((mul_34_17_n_7101 & mul_34_17_n_7102)
    | (mul_34_17_n_7102 & mul_34_17_n_7154)));
 assign mul_34_17_n_8148 = ((mul_34_17_n_7080 & mul_34_17_n_11494) | ((mul_34_17_n_7080 & mul_34_17_n_7084)
    | (mul_34_17_n_7084 & mul_34_17_n_11494)));
 assign mul_34_17_n_8146 = ((mul_34_17_n_6987 & mul_34_17_n_6356) | (mul_34_17_n_7634 & mul_34_17_n_5831));
 assign mul_34_17_n_8145 = ((mul_34_17_n_7098 & mul_34_17_n_7136) | ((mul_34_17_n_7098 & mul_34_17_n_5934)
    | (mul_34_17_n_5934 & mul_34_17_n_7136)));
 assign mul_34_17_n_8144 = ((mul_34_17_n_7114 & mul_34_17_n_6920) | ((mul_34_17_n_7114 & mul_34_17_n_22)
    | (mul_34_17_n_22 & mul_34_17_n_6920)));
 assign mul_34_17_n_8143 = ((mul_34_17_n_7073 & mul_34_17_n_7124) | ((mul_34_17_n_7073 & mul_34_17_n_110)
    | (mul_34_17_n_110 & mul_34_17_n_7124)));
 assign mul_34_17_n_8142 = ((mul_34_17_n_7297 & mul_34_17_n_6918) | ((mul_34_17_n_7297 & mul_34_17_n_6528)
    | (mul_34_17_n_6528 & mul_34_17_n_6918)));
 assign mul_34_17_n_8141 = ((mul_34_17_n_387 & mul_34_17_n_6631) | (mul_34_17_n_7613 & mul_34_17_n_5830));
 assign mul_34_17_n_8140 = ~(mul_34_17_n_7399 ^ mul_34_17_n_7142);
 assign mul_34_17_n_8138 = ~(mul_34_17_n_7400 ^ mul_34_17_n_7114);
 assign mul_34_17_n_8137 = (mul_34_17_n_7489 ^ mul_34_17_n_7794);
 assign mul_34_17_n_8136 = ((mul_34_17_n_196 & mul_34_17_n_7138) | ((mul_34_17_n_196 & mul_34_17_n_7298)
    | (mul_34_17_n_7298 & mul_34_17_n_7138)));
 assign mul_34_17_n_8135 = (mul_34_17_n_7468 ^ mul_34_17_n_7588);
 assign mul_34_17_n_8134 = (mul_34_17_n_7513 ^ mul_34_17_n_6779);
 assign mul_34_17_n_8133 = (mul_34_17_n_7572 ^ mul_34_17_n_191);
 assign mul_34_17_n_8132 = (mul_34_17_n_6787 ^ mul_34_17_n_7539);
 assign mul_34_17_n_8131 = ~((mul_34_17_n_7240 & mul_34_17_n_6355) | (mul_34_17_n_7640 & mul_34_17_n_5843));
 assign mul_34_17_n_8130 = ((mul_34_17_n_376 & mul_34_17_n_152) | (mul_34_17_n_7404 & mul_34_17_n_5828));
 assign mul_34_17_n_8129 = ((mul_34_17_n_7083 & mul_34_17_n_7144) | ((mul_34_17_n_7083 & mul_34_17_n_6900)
    | (mul_34_17_n_6900 & mul_34_17_n_7144)));
 assign mul_34_17_n_8127 = ~(mul_34_17_n_7402 ^ mul_34_17_n_7133);
 assign mul_34_17_n_8126 = ~((mul_34_17_n_6994 & mul_34_17_n_6354) | (mul_34_17_n_7641 & mul_34_17_n_5848));
 assign mul_34_17_n_8071 = ~mul_34_17_n_207;
 assign mul_34_17_n_8065 = ~mul_34_17_n_8064;
 assign mul_34_17_n_8054 = ~mul_34_17_n_8053;
 assign mul_34_17_n_8051 = ~mul_34_17_n_201;
 assign mul_34_17_n_8033 = ~mul_34_17_n_221;
 assign mul_34_17_n_8026 = ~mul_34_17_n_8027;
 assign mul_34_17_n_8021 = ~mul_34_17_n_8020;
 assign mul_34_17_n_8005 = ~mul_34_17_n_8004;
 assign mul_34_17_n_7993 = ~mul_34_17_n_218;
 assign mul_34_17_n_7987 = ~mul_34_17_n_164;
 assign mul_34_17_n_7979 = ~mul_34_17_n_7980;
 assign mul_34_17_n_7978 = ~(mul_34_17_n_7414 | mul_34_17_n_7684);
 assign mul_34_17_n_7976 = ~(mul_34_17_n_7079 ^ mul_34_17_n_7310);
 assign mul_34_17_n_7975 = ~(mul_34_17_n_7159 ^ mul_34_17_n_6404);
 assign mul_34_17_n_7974 = ((mul_34_17_n_6403 & mul_34_17_n_7384) | ((mul_34_17_n_6403 & mul_34_17_n_5465)
    | (mul_34_17_n_5465 & mul_34_17_n_7384)));
 assign mul_34_17_n_7973 = ~(mul_34_17_n_7768 | mul_34_17_n_6921);
 assign mul_34_17_n_7972 = ~((mul_34_17_n_7286 & mul_34_17_n_7287) | (mul_34_17_n_7389 & mul_34_17_n_7252));
 assign mul_34_17_n_7971 = ~(mul_34_17_n_7589 | mul_34_17_n_7596);
 assign mul_34_17_n_7970 = ~(mul_34_17_n_7598 | mul_34_17_n_6776);
 assign mul_34_17_n_7968 = (mul_34_17_n_7079 ^ mul_34_17_n_7310);
 assign mul_34_17_n_7964 = ~(mul_34_17_n_7064 ^ mul_34_17_n_7055);
 assign mul_34_17_n_7963 = ~(mul_34_17_n_194 ^ mul_34_17_n_6492);
 assign mul_34_17_n_7961 = ~(mul_34_17_n_7321 ^ mul_34_17_n_5983);
 assign mul_34_17_n_7960 = ~(mul_34_17_n_7326 ^ mul_34_17_n_7341);
 assign mul_34_17_n_7959 = ~(mul_34_17_n_7414 & mul_34_17_n_7684);
 assign mul_34_17_n_7958 = (mul_34_17_n_7078 ^ mul_34_17_n_6794);
 assign mul_34_17_n_7957 = (mul_34_17_n_196 ^ mul_34_17_n_7298);
 assign mul_34_17_n_7956 = (mul_34_17_n_176 ^ mul_34_17_n_7362);
 assign mul_34_17_n_7955 = (mul_34_17_n_7323 ^ mul_34_17_n_7324);
 assign mul_34_17_n_7954 = ~(mul_34_17_n_7358 ^ mul_34_17_n_7334);
 assign mul_34_17_n_7953 = (mul_34_17_n_6778 ^ mul_34_17_n_7359);
 assign mul_34_17_n_8072 = ((mul_34_17_n_6407 & mul_34_17_n_6686) | (mul_34_17_n_7159 & mul_34_17_n_6404));
 assign mul_34_17_n_7952 = (mul_34_17_n_7355 ^ mul_34_17_n_7332);
 assign mul_34_17_n_8070 = ~((mul_34_17_n_6307 | mul_34_17_n_5987) & (mul_34_17_n_7164 | mul_34_17_n_6933));
 assign mul_34_17_n_8069 = (mul_34_17_n_7153 ^ mul_34_17_n_7322);
 assign mul_34_17_n_7951 = (mul_34_17_n_198 ^ mul_34_17_n_7307);
 assign mul_34_17_n_7950 = ~(mul_34_17_n_7149 ^ mul_34_17_n_6911);
 assign mul_34_17_n_7949 = ~(mul_34_17_n_7293 ^ mul_34_17_n_6476);
 assign mul_34_17_n_7948 = (mul_34_17_n_7144 ^ mul_34_17_n_6900);
 assign mul_34_17_n_7947 = (mul_34_17_n_7377 ^ mul_34_17_n_6901);
 assign mul_34_17_n_8068 = ~(mul_34_17_n_7802 & mul_34_17_n_7365);
 assign mul_34_17_n_8067 = ((mul_34_17_n_6931 & mul_34_17_n_6814) | ((mul_34_17_n_6931 & mul_34_17_n_5202)
    | (mul_34_17_n_5202 & mul_34_17_n_6814)));
 assign mul_34_17_n_8066 = ~(mul_34_17_n_7074 ^ mul_34_17_n_6176);
 assign mul_34_17_n_7946 = (mul_34_17_n_7328 ^ mul_34_17_n_6575);
 assign mul_34_17_n_8064 = ~(mul_34_17_n_6547 ^ (mul_34_17_n_6670 ^ (mul_34_17_n_5487 ^ mul_34_17_n_4401)));
 assign mul_34_17_n_8063 = ((mul_34_17_n_6891 & mul_34_17_n_6679) | (mul_34_17_n_7285 & mul_34_17_n_5814));
 assign mul_34_17_n_8062 = ((mul_34_17_n_6605 & mul_34_17_n_7344) | ((mul_34_17_n_6605 & mul_34_17_n_6904)
    | (mul_34_17_n_6904 & mul_34_17_n_7344)));
 assign mul_34_17_n_8061 = ((mul_34_17_n_6890 & mul_34_17_n_6688) | (mul_34_17_n_7281 & mul_34_17_n_5858));
 assign mul_34_17_n_8060 = ((mul_34_17_n_6884 | mul_34_17_n_147) & (mul_34_17_n_7268 | mul_34_17_n_5851));
 assign mul_34_17_n_8059 = ((mul_34_17_n_7 & mul_34_17_n_7148) | ((mul_34_17_n_7 & mul_34_17_n_5708)
    | (mul_34_17_n_5708 & mul_34_17_n_7148)));
 assign mul_34_17_n_8057 = ~(mul_34_17_n_6936 ^ mul_34_17_n_6162);
 assign mul_34_17_n_8056 = ~(mul_34_17_n_7089 ^ mul_34_17_n_102);
 assign mul_34_17_n_8055 = ~(mul_34_17_n_7081 ^ mul_34_17_n_119);
 assign mul_34_17_n_8053 = ~(mul_34_17_n_7314 ^ mul_34_17_n_6520);
 assign mul_34_17_n_8052 = ~((mul_34_17_n_7046 & ~mul_34_17_n_6664) | (mul_34_17_n_7265 & mul_34_17_n_6664));
 assign mul_34_17_n_8050 = ((mul_34_17_n_6915 & mul_34_17_n_194) | ((mul_34_17_n_6915 & mul_34_17_n_6491)
    | (mul_34_17_n_6491 & mul_34_17_n_194)));
 assign mul_34_17_n_8049 = ~(mul_34_17_n_6639 ^ (mul_34_17_n_6600 ^ (mul_34_17_n_5474 ^ mul_34_17_n_4753)));
 assign mul_34_17_n_8048 = ~(mul_34_17_n_7189 ^ mul_34_17_n_5798);
 assign mul_34_17_n_8046 = ~(mul_34_17_n_7169 ^ mul_34_17_n_6659);
 assign mul_34_17_n_8044 = ~(mul_34_17_n_7188 ^ mul_34_17_n_7343);
 assign mul_34_17_n_8042 = ((mul_34_17_n_389 & mul_34_17_n_6636) | (mul_34_17_n_7283 & mul_34_17_n_5861));
 assign mul_34_17_n_8041 = (mul_34_17_n_6909 ^ mul_34_17_n_7370);
 assign mul_34_17_n_8040 = ((mul_34_17_n_6611 & mul_34_17_n_7361) | ((mul_34_17_n_6611 & mul_34_17_n_5551)
    | (mul_34_17_n_5551 & mul_34_17_n_7361)));
 assign mul_34_17_n_8037 = (mul_34_17_n_7375 ^ mul_34_17_n_7295);
 assign mul_34_17_n_8036 = ((mul_34_17_n_6786 & mul_34_17_n_7155) | ((mul_34_17_n_6786 & mul_34_17_n_5968)
    | (mul_34_17_n_5968 & mul_34_17_n_7155)));
 assign mul_34_17_n_8035 = ~(mul_34_17_n_7174 ^ mul_34_17_n_5704);
 assign mul_34_17_n_8032 = ~(mul_34_17_n_7171 ^ mul_34_17_n_6922);
 assign mul_34_17_n_8031 = ~(mul_34_17_n_7170 ^ mul_34_17_n_5698);
 assign mul_34_17_n_8030 = ((mul_34_17_n_6253 & mul_34_17_n_7134) | ((mul_34_17_n_6253 & mul_34_17_n_6784)
    | (mul_34_17_n_6784 & mul_34_17_n_7134)));
 assign mul_34_17_n_8028 = ((mul_34_17_n_6134 & mul_34_17_n_7372) | ((mul_34_17_n_6134 & mul_34_17_n_6137)
    | (mul_34_17_n_6137 & mul_34_17_n_7372)));
 assign mul_34_17_n_8027 = ~(mul_34_17_n_7347 ^ mul_34_17_n_5944);
 assign mul_34_17_n_8025 = ~(mul_34_17_n_7166 ^ mul_34_17_n_5769);
 assign mul_34_17_n_8024 = ~(mul_34_17_n_6943 ^ mul_34_17_n_5988);
 assign mul_34_17_n_8023 = ((mul_34_17_n_6417 & mul_34_17_n_7151) | ((mul_34_17_n_6417 & mul_34_17_n_6418)
    | (mul_34_17_n_6418 & mul_34_17_n_7151)));
 assign mul_34_17_n_8022 = ~(mul_34_17_n_7173 ^ mul_34_17_n_6919);
 assign mul_34_17_n_8020 = ((mul_34_17_n_37 & mul_34_17_n_7147) | ((mul_34_17_n_37 & mul_34_17_n_6277)
    | (mul_34_17_n_6277 & mul_34_17_n_7147)));
 assign mul_34_17_n_8019 = ~(mul_34_17_n_7175 ^ mul_34_17_n_5677);
 assign mul_34_17_n_8017 = ~(mul_34_17_n_151 ^ mul_34_17_n_108);
 assign mul_34_17_n_8016 = ~(mul_34_17_n_6948 ^ mul_34_17_n_5630);
 assign mul_34_17_n_8015 = ((mul_34_17_n_7284 & mul_34_17_n_72) | (mul_34_17_n_7266 & mul_34_17_n_6683));
 assign mul_34_17_n_8013 = ((mul_34_17_n_6897 & mul_34_17_n_7345) | ((mul_34_17_n_6897 & mul_34_17_n_6566)
    | (mul_34_17_n_6566 & mul_34_17_n_7345)));
 assign mul_34_17_n_8012 = ((mul_34_17_n_7020 & mul_34_17_n_6406) | (mul_34_17_n_7246 & mul_34_17_n_6405));
 assign mul_34_17_n_8011 = (mul_34_17_n_7301 ^ mul_34_17_n_7364);
 assign mul_34_17_n_8010 = ~(mul_34_17_n_7179 ^ mul_34_17_n_7150);
 assign mul_34_17_n_8009 = ((mul_34_17_n_11514 & mul_34_17_n_7342) | ((mul_34_17_n_11514 & mul_34_17_n_1)
    | (mul_34_17_n_1 & mul_34_17_n_7342)));
 assign mul_34_17_n_8008 = ((mul_34_17_n_6789 & mul_34_17_n_7291) | ((mul_34_17_n_6789 & mul_34_17_n_6497)
    | (mul_34_17_n_6497 & mul_34_17_n_7291)));
 assign mul_34_17_n_8007 = ~(mul_34_17_n_6947 ^ mul_34_17_n_6391);
 assign mul_34_17_n_8004 = ((mul_34_17_n_84 & mul_34_17_n_7139) | ((mul_34_17_n_84 & mul_34_17_n_83)
    | (mul_34_17_n_83 & mul_34_17_n_7139)));
 assign mul_34_17_n_8003 = ~(mul_34_17_n_7167 ^ mul_34_17_n_5668);
 assign mul_34_17_n_8002 = ~(mul_34_17_n_7387 ^ mul_34_17_n_5649);
 assign mul_34_17_n_8001 = (mul_34_17_n_7320 ^ mul_34_17_n_6649);
 assign mul_34_17_n_7998 = ~(mul_34_17_n_7177 ^ mul_34_17_n_6629);
 assign mul_34_17_n_7996 = ((mul_34_17_n_6673 & mul_34_17_n_7343) | ((mul_34_17_n_6673 & mul_34_17_n_94)
    | (mul_34_17_n_94 & mul_34_17_n_7343)));
 assign mul_34_17_n_7986 = ~(mul_34_17_n_6938 ^ mul_34_17_n_5710);
 assign mul_34_17_n_7984 = ~((mul_34_17_n_7199 & ~mul_34_17_n_6349) | (mul_34_17_n_7242 & mul_34_17_n_6349));
 assign mul_34_17_n_7983 = (mul_34_17_n_7386 ^ mul_34_17_n_5912);
 assign mul_34_17_n_7981 = ~((mul_34_17_n_7019 & ~mul_34_17_n_6392) | (mul_34_17_n_7259 & mul_34_17_n_6392));
 assign mul_34_17_n_7980 = ~(mul_34_17_n_6949 ^ mul_34_17_n_7152);
 assign mul_34_17_n_7944 = ~mul_34_17_n_7943;
 assign mul_34_17_n_7931 = ~mul_34_17_n_7930;
 assign mul_34_17_n_7928 = ~mul_34_17_n_7927;
 assign mul_34_17_n_7925 = ~mul_34_17_n_7924;
 assign mul_34_17_n_7923 = ~mul_34_17_n_206;
 assign mul_34_17_n_7918 = ~mul_34_17_n_7919;
 assign mul_34_17_n_7915 = ~mul_34_17_n_11428;
 assign mul_34_17_n_7901 = ~mul_34_17_n_7902;
 assign mul_34_17_n_7897 = ~mul_34_17_n_7896;
 assign mul_34_17_n_7890 = ~mul_34_17_n_7889;
 assign mul_34_17_n_7878 = ~mul_34_17_n_7877;
 assign mul_34_17_n_7862 = ~mul_34_17_n_7861;
 assign mul_34_17_n_7857 = ~mul_34_17_n_7858;
 assign mul_34_17_n_7844 = ~mul_34_17_n_7843;
 assign mul_34_17_n_7836 = ~mul_34_17_n_180;
 assign mul_34_17_n_7834 = ~mul_34_17_n_7835;
 assign mul_34_17_n_7824 = (mul_34_17_n_7052 ^ mul_34_17_n_7059);
 assign mul_34_17_n_7823 = ~(mul_34_17_n_7059 ^ mul_34_17_n_7052);
 assign mul_34_17_n_7821 = (mul_34_17_n_187 ^ mul_34_17_n_6914);
 assign mul_34_17_n_7820 = (mul_34_17_n_7304 ^ mul_34_17_n_6802);
 assign mul_34_17_n_7819 = (mul_34_17_n_7124 ^ mul_34_17_n_110);
 assign mul_34_17_n_7945 = ~(mul_34_17_n_7086 ^ mul_34_17_n_7062);
 assign mul_34_17_n_7943 = ~(mul_34_17_n_7088 ^ mul_34_17_n_6175);
 assign mul_34_17_n_7942 = (mul_34_17_n_7105 ^ mul_34_17_n_6331);
 assign mul_34_17_n_7818 = ~(mul_34_17_n_7382 ^ mul_34_17_n_6780);
 assign mul_34_17_n_7941 = ~(mul_34_17_n_7342 ^ mul_34_17_n_7184);
 assign mul_34_17_n_7817 = (mul_34_17_n_5934 ^ mul_34_17_n_7136);
 assign mul_34_17_n_7816 = (mul_34_17_n_7135 ^ mul_34_17_n_5707);
 assign mul_34_17_n_7815 = (mul_34_17_n_7125 ^ mul_34_17_n_7099);
 assign mul_34_17_n_7814 = (mul_34_17_n_7367 ^ mul_34_17_n_7333);
 assign mul_34_17_n_7940 = (mul_34_17_n_7154 ^ mul_34_17_n_7101);
 assign mul_34_17_n_7939 = (mul_34_17_n_7374 ^ mul_34_17_n_7352);
 assign mul_34_17_n_7938 = ~(mul_34_17_n_5987 ^ (mul_34_17_n_6307 ^ (mul_34_17_n_6309 ^ mul_34_17_n_5108)));
 assign mul_34_17_n_7813 = ~(mul_34_17_n_7126 ^ mul_34_17_n_59);
 assign mul_34_17_n_7937 = ~(mul_34_17_n_7108 ^ mul_34_17_n_6508);
 assign mul_34_17_n_7812 = (mul_34_17_n_199 ^ mul_34_17_n_171);
 assign mul_34_17_n_7811 = (mul_34_17_n_7338 ^ mul_34_17_n_11520);
 assign mul_34_17_n_7810 = (mul_34_17_n_7120 ^ mul_34_17_n_7077);
 assign mul_34_17_n_7809 = (mul_34_17_n_7080 ^ mul_34_17_n_7084);
 assign mul_34_17_n_7936 = (mul_34_17_n_11643 ^ mul_34_17_n_7327);
 assign mul_34_17_n_7808 = (mul_34_17_n_7308 ^ mul_34_17_n_6616);
 assign mul_34_17_n_7935 = ~((mul_34_17_n_7000 & ~mul_34_17_n_6251) | (mul_34_17_n_6995 & mul_34_17_n_6251));
 assign mul_34_17_n_7934 = ~(mul_34_17_n_7104 ^ mul_34_17_n_6490);
 assign mul_34_17_n_7933 = ~(mul_34_17_n_7093 ^ mul_34_17_n_6173);
 assign mul_34_17_n_7932 = ~(mul_34_17_n_6966 ^ mul_34_17_n_123);
 assign mul_34_17_n_7930 = ~(mul_34_17_n_7110 ^ mul_34_17_n_6194);
 assign mul_34_17_n_7929 = ~(mul_34_17_n_7112 ^ mul_34_17_n_55);
 assign mul_34_17_n_7927 = ~(mul_34_17_n_7117 ^ mul_34_17_n_6186);
 assign mul_34_17_n_7807 = ~(mul_34_17_n_6394 ^ (mul_34_17_n_6246 ^ (mul_34_17_n_5153 ^ mul_34_17_n_3764)));
 assign mul_34_17_n_7806 = (mul_34_17_n_7158 ^ mul_34_17_n_5530);
 assign mul_34_17_n_7926 = ((mul_34_17_n_6234 & mul_34_17_n_7063) | ((mul_34_17_n_6234 & mul_34_17_n_5705)
    | (mul_34_17_n_5705 & mul_34_17_n_7063)));
 assign mul_34_17_n_7924 = ~(mul_34_17_n_6302 ^ (mul_34_17_n_6303 ^ (mul_34_17_n_5193 ^ mul_34_17_n_4699)));
 assign mul_34_17_n_7922 = ~((mul_34_17_n_7194 & ~mul_34_17_n_6567) | (mul_34_17_n_7193 & mul_34_17_n_6567));
 assign mul_34_17_n_7919 = ~(mul_34_17_n_6951 ^ mul_34_17_n_6917);
 assign mul_34_17_n_7913 = ~((mul_34_17_n_6974 & ~mul_34_17_n_6577) | (mul_34_17_n_7288 & mul_34_17_n_6577));
 assign mul_34_17_n_7911 = ~((mul_34_17_n_6171 & (~mul_34_17_n_6212 & ~mul_34_17_n_6231)) | ((mul_34_17_n_6170
    & (mul_34_17_n_6212 & ~mul_34_17_n_6231)) | (mul_34_17_n_7022 & mul_34_17_n_6231)));
 assign mul_34_17_n_7908 = ~((mul_34_17_n_5411 & (~mul_34_17_n_6198 & ~mul_34_17_n_6297)) | ((mul_34_17_n_5410
    & (mul_34_17_n_6198 & ~mul_34_17_n_6297)) | (mul_34_17_n_7012 & mul_34_17_n_6297)));
 assign mul_34_17_n_7906 = ~((mul_34_17_n_136 & (~mul_34_17_n_6504 & ~mul_34_17_n_6562)) | ((mul_34_17_n_6493
    & (mul_34_17_n_6504 & ~mul_34_17_n_6562)) | (mul_34_17_n_7002 & mul_34_17_n_6562)));
 assign mul_34_17_n_7905 = ~((mul_34_17_n_6978 & ~mul_34_17_n_6327) | (mul_34_17_n_6979 & mul_34_17_n_6327));
 assign mul_34_17_n_7903 = ~((mul_34_17_n_7255 & ~mul_34_17_n_6352) | (mul_34_17_n_7024 & mul_34_17_n_6352));
 assign mul_34_17_n_7902 = ~(mul_34_17_n_6950 ^ mul_34_17_n_5897);
 assign mul_34_17_n_7900 = ~(mul_34_17_n_6960 ^ mul_34_17_n_5568);
 assign mul_34_17_n_7899 = ((mul_34_17_n_6260 & mul_34_17_n_7131) | ((mul_34_17_n_6260 & mul_34_17_n_21)
    | (mul_34_17_n_21 & mul_34_17_n_7131)));
 assign mul_34_17_n_7898 = ((mul_34_17_n_6615 & mul_34_17_n_7360) | ((mul_34_17_n_6615 & mul_34_17_n_6905)
    | (mul_34_17_n_6905 & mul_34_17_n_7360)));
 assign mul_34_17_n_7896 = ~((mul_34_17_n_3986 & (~mul_34_17_n_5418 & ~mul_34_17_n_7187)) | ((mul_34_17_n_3985
    & (mul_34_17_n_5418 & ~mul_34_17_n_7187)) | (mul_34_17_n_6647 & mul_34_17_n_7187)));
 assign mul_34_17_n_7895 = ~((mul_34_17_n_6595 & (~mul_34_17_n_5427 & ~mul_34_17_n_7185)) | ((mul_34_17_n_6596
    & (mul_34_17_n_5427 & ~mul_34_17_n_7185)) | (mul_34_17_n_7198 & mul_34_17_n_7185)));
 assign mul_34_17_n_7894 = ((mul_34_17_n_6236 & mul_34_17_n_7152) | ((mul_34_17_n_6236 & mul_34_17_n_5714)
    | (mul_34_17_n_5714 & mul_34_17_n_7152)));
 assign mul_34_17_n_7893 = ~((mul_34_17_n_5432 & (~mul_34_17_n_3982 & ~mul_34_17_n_6937)) | ((mul_34_17_n_5433
    & (mul_34_17_n_3982 & ~mul_34_17_n_6937)) | (mul_34_17_n_6654 & mul_34_17_n_6937)));
 assign mul_34_17_n_7889 = ((mul_34_17_n_6532 & mul_34_17_n_7142) | ((mul_34_17_n_6532 & mul_34_17_n_6777)
    | (mul_34_17_n_6777 & mul_34_17_n_7142)));
 assign mul_34_17_n_7888 = ((mul_34_17_n_6318 & mul_34_17_n_174) | ((mul_34_17_n_6318 & mul_34_17_n_5595)
    | (mul_34_17_n_5595 & mul_34_17_n_174)));
 assign mul_34_17_n_7887 = ~(mul_34_17_n_7388 ^ mul_34_17_n_6074);
 assign mul_34_17_n_7885 = ~(mul_34_17_n_7804 & mul_34_17_n_6935);
 assign mul_34_17_n_7884 = ~((mul_34_17_n_7256 & ~mul_34_17_n_6350) | (mul_34_17_n_6985 & mul_34_17_n_6350));
 assign mul_34_17_n_7882 = ~(mul_34_17_n_6965 ^ mul_34_17_n_6797);
 assign mul_34_17_n_7881 = ~((mul_34_17_n_7218 & ~mul_34_17_n_6597) | (mul_34_17_n_7217 & mul_34_17_n_6597));
 assign mul_34_17_n_7880 = ~(mul_34_17_n_6963 ^ mul_34_17_n_7372);
 assign mul_34_17_n_7877 = ~(mul_34_17_n_6962 ^ mul_34_17_n_174);
 assign mul_34_17_n_7876 = ((mul_34_17_n_6241 & mul_34_17_n_7141) | ((mul_34_17_n_6241 & mul_34_17_n_6242)
    | (mul_34_17_n_6242 & mul_34_17_n_7141)));
 assign mul_34_17_n_7875 = ~((mul_34_17_n_7237 & ~mul_34_17_n_6542) | (mul_34_17_n_7233 & mul_34_17_n_6542));
 assign mul_34_17_n_7872 = ~(mul_34_17_n_6955 ^ mul_34_17_n_7130);
 assign mul_34_17_n_7871 = ~(mul_34_17_n_6956 ^ mul_34_17_n_5116);
 assign mul_34_17_n_7869 = ~(mul_34_17_n_6964 ^ mul_34_17_n_5531);
 assign mul_34_17_n_7867 = ~(mul_34_17_n_6959 ^ mul_34_17_n_73);
 assign mul_34_17_n_7865 = ~(mul_34_17_n_6946 ^ mul_34_17_n_6641);
 assign mul_34_17_n_7864 = ~(mul_34_17_n_6957 ^ mul_34_17_n_5922);
 assign mul_34_17_n_7861 = ~(mul_34_17_n_7092 ^ mul_34_17_n_7072);
 assign mul_34_17_n_7860 = ~(mul_34_17_n_6954 ^ mul_34_17_n_7147);
 assign mul_34_17_n_7805 = ~(mul_34_17_n_7157 ^ mul_34_17_n_5719);
 assign mul_34_17_n_7858 = ((mul_34_17_n_6323 & mul_34_17_n_7132) | ((mul_34_17_n_6323 & mul_34_17_n_6239)
    | (mul_34_17_n_6239 & mul_34_17_n_7132)));
 assign mul_34_17_n_7855 = ~((mul_34_17_n_6188 & mul_34_17_n_6295) | (mul_34_17_n_6971 & mul_34_17_n_5834));
 assign mul_34_17_n_7854 = ~((mul_34_17_n_6487 & (~mul_34_17_n_6517 & ~mul_34_17_n_6573)) | ((mul_34_17_n_6486
    & (mul_34_17_n_6517 & ~mul_34_17_n_6573)) | (mul_34_17_n_6975 & mul_34_17_n_6573)));
 assign mul_34_17_n_7853 = ~((mul_34_17_n_7249 & ~mul_34_17_n_6387) | (mul_34_17_n_6983 & mul_34_17_n_6387));
 assign mul_34_17_n_7852 = ~((mul_34_17_n_7011 & ~mul_34_17_n_6268) | (mul_34_17_n_7014 & mul_34_17_n_6268));
 assign mul_34_17_n_7850 = ~((mul_34_17_n_145 & (~mul_34_17_n_6511 & ~mul_34_17_n_6531)) | ((mul_34_17_n_6455
    & (mul_34_17_n_6511 & ~mul_34_17_n_6531)) | (mul_34_17_n_7195 & mul_34_17_n_6531)));
 assign mul_34_17_n_7846 = ~((mul_34_17_n_7282 & ~mul_34_17_n_6626) | (mul_34_17_n_7207 & mul_34_17_n_6626));
 assign mul_34_17_n_7845 = ~((mul_34_17_n_6989 & ~mul_34_17_n_6317) | (mul_34_17_n_6990 & mul_34_17_n_6317));
 assign mul_34_17_n_7843 = ~((mul_34_17_n_7048 & ~mul_34_17_n_6223) | (mul_34_17_n_7043 & mul_34_17_n_6223));
 assign mul_34_17_n_7842 = ~((mul_34_17_n_5413 & (~mul_34_17_n_6524 & ~mul_34_17_n_6576)) | ((mul_34_17_n_5412
    & (mul_34_17_n_6524 & ~mul_34_17_n_6576)) | (mul_34_17_n_7220 & mul_34_17_n_6576)));
 assign mul_34_17_n_7839 = ~((mul_34_17_n_5423 & (~mul_34_17_n_3072 & ~mul_34_17_n_7183)) | ((mul_34_17_n_5424
    & (mul_34_17_n_3072 & ~mul_34_17_n_7183)) | (mul_34_17_n_6634 & mul_34_17_n_7183)));
 assign mul_34_17_n_7838 = ~((mul_34_17_n_3065 & (~mul_34_17_n_5121 & ~mul_34_17_n_7186)) | ((mul_34_17_n_3066
    & (mul_34_17_n_5121 & ~mul_34_17_n_7186)) | (mul_34_17_n_6395 & mul_34_17_n_7186)));
 assign mul_34_17_n_7835 = ~(mul_34_17_n_6945 ^ mul_34_17_n_5706);
 assign mul_34_17_n_7832 = ~(mul_34_17_n_6961 ^ mul_34_17_n_43);
 assign mul_34_17_n_7803 = ~mul_34_17_n_7802;
 assign mul_34_17_n_7780 = ~mul_34_17_n_7781;
 assign mul_34_17_n_7774 = ~mul_34_17_n_7773;
 assign mul_34_17_n_7755 = ~mul_34_17_n_7754;
 assign mul_34_17_n_7753 = ~mul_34_17_n_162;
 assign mul_34_17_n_7750 = ~mul_34_17_n_7751;
 assign mul_34_17_n_7745 = ~mul_34_17_n_7744;
 assign mul_34_17_n_7729 = ~mul_34_17_n_7728;
 assign mul_34_17_n_7721 = ~mul_34_17_n_7720;
 assign mul_34_17_n_7718 = ~mul_34_17_n_7717;
 assign mul_34_17_n_7709 = ~mul_34_17_n_7708;
 assign mul_34_17_n_7681 = ~mul_34_17_n_7680;
 assign mul_34_17_n_7675 = ~mul_34_17_n_7674;
 assign mul_34_17_n_7672 = ~mul_34_17_n_7673;
 assign mul_34_17_n_7665 = ~(mul_34_17_n_383 | mul_34_17_n_5862);
 assign mul_34_17_n_7664 = ~(mul_34_17_n_7303 | mul_34_17_n_6457);
 assign mul_34_17_n_7663 = ~(mul_34_17_n_7303 & mul_34_17_n_6457);
 assign mul_34_17_n_7662 = ~(mul_34_17_n_7210 | mul_34_17_n_5859);
 assign mul_34_17_n_7661 = ~(mul_34_17_n_7305 & mul_34_17_n_6477);
 assign mul_34_17_n_7660 = ~(mul_34_17_n_7374 & mul_34_17_n_7352);
 assign mul_34_17_n_7659 = ~(mul_34_17_n_7296 & mul_34_17_n_6465);
 assign mul_34_17_n_7658 = ~(mul_34_17_n_7296 | mul_34_17_n_6465);
 assign mul_34_17_n_7657 = ~(mul_34_17_n_7111 | mul_34_17_n_26);
 assign mul_34_17_n_7656 = ~(mul_34_17_n_381 | mul_34_17_n_5854);
 assign mul_34_17_n_7655 = ~(mul_34_17_n_382 | mul_34_17_n_5852);
 assign mul_34_17_n_7654 = ~(mul_34_17_n_7314 & mul_34_17_n_6519);
 assign mul_34_17_n_7653 = ~(mul_34_17_n_7314 | mul_34_17_n_6519);
 assign mul_34_17_n_7652 = ~(mul_34_17_n_7244 | mul_34_17_n_6443);
 assign mul_34_17_n_7651 = ~(mul_34_17_n_7089 & mul_34_17_n_102);
 assign mul_34_17_n_7650 = ~(mul_34_17_n_7089 | mul_34_17_n_102);
 assign mul_34_17_n_7649 = ~(mul_34_17_n_7081 | mul_34_17_n_119);
 assign mul_34_17_n_7648 = ~(mul_34_17_n_7081 & mul_34_17_n_119);
 assign mul_34_17_n_7647 = ~(mul_34_17_n_7027 | mul_34_17_n_5847);
 assign mul_34_17_n_7646 = ~(mul_34_17_n_7094 & mul_34_17_n_6161);
 assign mul_34_17_n_7645 = ~(mul_34_17_n_7094 | mul_34_17_n_6161);
 assign mul_34_17_n_7644 = ~(mul_34_17_n_6970 | mul_34_17_n_6124);
 assign mul_34_17_n_7643 = ~(mul_34_17_n_7067 | mul_34_17_n_6200);
 assign mul_34_17_n_7642 = ~(mul_34_17_n_379 | mul_34_17_n_6121);
 assign mul_34_17_n_7641 = ~(mul_34_17_n_6993 | mul_34_17_n_5849);
 assign mul_34_17_n_7640 = ~(mul_34_17_n_6992 | mul_34_17_n_5842);
 assign mul_34_17_n_7639 = ~(mul_34_17_n_7112 & mul_34_17_n_55);
 assign mul_34_17_n_7638 = ~(mul_34_17_n_7112 | mul_34_17_n_55);
 assign mul_34_17_n_7637 = ~(mul_34_17_n_7117 & mul_34_17_n_6185);
 assign mul_34_17_n_7636 = ~(mul_34_17_n_7110 & mul_34_17_n_6193);
 assign mul_34_17_n_7635 = ~(mul_34_17_n_7111 & mul_34_17_n_26);
 assign mul_34_17_n_7634 = ~(mul_34_17_n_6969 | mul_34_17_n_5841);
 assign mul_34_17_n_7633 = ~(mul_34_17_n_7110 | mul_34_17_n_6193);
 assign mul_34_17_n_7804 = ~(mul_34_17_n_6984 & mul_34_17_n_4884);
 assign mul_34_17_n_7632 = ~(mul_34_17_n_7388 & mul_34_17_n_6074);
 assign mul_34_17_n_7631 = ~(mul_34_17_n_6854 & (mul_34_17_n_6826 & (mul_34_17_n_5500 & mul_34_17_n_4904)));
 assign mul_34_17_n_7630 = ~(mul_34_17_n_7208 | mul_34_17_n_6447);
 assign mul_34_17_n_7629 = ~(mul_34_17_n_385 | mul_34_17_n_6441);
 assign mul_34_17_n_7628 = ~(mul_34_17_n_7190 | mul_34_17_n_5866);
 assign mul_34_17_n_7627 = ~(mul_34_17_n_7162 & mul_34_17_n_7161);
 assign mul_34_17_n_7626 = ~(mul_34_17_n_7117 | mul_34_17_n_6185);
 assign mul_34_17_n_7625 = ~(mul_34_17_n_7163 & mul_34_17_n_7160);
 assign mul_34_17_n_7624 = ~(mul_34_17_n_6931 ^ mul_34_17_n_5202);
 assign mul_34_17_n_7623 = ~((mul_34_17_n_6184 | mul_34_17_n_6177) & (mul_34_17_n_6832 | mul_34_17_n_6405));
 assign mul_34_17_n_7622 = ~(mul_34_17_n_7164 | mul_34_17_n_6933);
 assign mul_34_17_n_7621 = ~(mul_34_17_n_7108 & mul_34_17_n_6508);
 assign mul_34_17_n_7620 = ~(mul_34_17_n_7108 | mul_34_17_n_6508);
 assign mul_34_17_n_7619 = ~(mul_34_17_n_388 | mul_34_17_n_5835);
 assign mul_34_17_n_7618 = ~(mul_34_17_n_6976 | mul_34_17_n_6434);
 assign mul_34_17_n_7617 = ~(mul_34_17_n_7104 & mul_34_17_n_6490);
 assign mul_34_17_n_7616 = ~(mul_34_17_n_7104 | mul_34_17_n_6490);
 assign mul_34_17_n_7615 = ~(mul_34_17_n_7093 & mul_34_17_n_6173);
 assign mul_34_17_n_7614 = ~(mul_34_17_n_7093 | mul_34_17_n_6173);
 assign mul_34_17_n_7613 = ~(mul_34_17_n_387 | mul_34_17_n_5829);
 assign mul_34_17_n_7612 = ~(mul_34_17_n_7086 & mul_34_17_n_7062);
 assign mul_34_17_n_7611 = ~(mul_34_17_n_7086 | mul_34_17_n_7062);
 assign mul_34_17_n_7610 = ~(mul_34_17_n_7067 & mul_34_17_n_6200);
 assign mul_34_17_n_7609 = ~(mul_34_17_n_7088 & mul_34_17_n_6175);
 assign mul_34_17_n_7608 = ~(mul_34_17_n_7088 | mul_34_17_n_6175);
 assign mul_34_17_n_7607 = ~(mul_34_17_n_7074 & mul_34_17_n_6176);
 assign mul_34_17_n_7606 = ~(mul_34_17_n_7074 | mul_34_17_n_6176);
 assign mul_34_17_n_7802 = ((mul_34_17_n_6403 | mul_34_17_n_5465) & (mul_34_17_n_6888 | mul_34_17_n_204));
 assign mul_34_17_n_7605 = (mul_34_17_n_6615 ^ mul_34_17_n_6905);
 assign mul_34_17_n_7801 = ((mul_34_17_n_6570 & mul_34_17_n_154) | ((mul_34_17_n_6570 & mul_34_17_n_6571)
    | (mul_34_17_n_6571 & mul_34_17_n_154)));
 assign mul_34_17_n_7604 = (mul_34_17_n_6605 ^ mul_34_17_n_6904);
 assign mul_34_17_n_7603 = ((mul_34_17_n_6458 & mul_34_17_n_6498) | ((mul_34_17_n_6458 & mul_34_17_n_6559)
    | (mul_34_17_n_6559 & mul_34_17_n_6498)));
 assign mul_34_17_n_7602 = ((mul_34_17_n_6459 & mul_34_17_n_6503) | ((mul_34_17_n_6459 & mul_34_17_n_6563)
    | (mul_34_17_n_6563 & mul_34_17_n_6503)));
 assign mul_34_17_n_7800 = ((mul_34_17_n_142 & mul_34_17_n_34) | ((mul_34_17_n_142 & mul_34_17_n_122)
    | (mul_34_17_n_122 & mul_34_17_n_34)));
 assign mul_34_17_n_7799 = ((mul_34_17_n_71 & mul_34_17_n_6502) | ((mul_34_17_n_71 & mul_34_17_n_6461)
    | (mul_34_17_n_6461 & mul_34_17_n_6502)));
 assign mul_34_17_n_7798 = ((mul_34_17_n_35 & mul_34_17_n_6797) | ((mul_34_17_n_35 & mul_34_17_n_36)
    | (mul_34_17_n_36 & mul_34_17_n_6797)));
 assign mul_34_17_n_7797 = ((mul_34_17_n_6560 & mul_34_17_n_6650) | ((mul_34_17_n_6560 & mul_34_17_n_5133)
    | (mul_34_17_n_5133 & mul_34_17_n_6650)));
 assign mul_34_17_n_7601 = ~(mul_34_17_n_7159 | mul_34_17_n_6404);
 assign mul_34_17_n_7796 = ((mul_34_17_n_6301 & mul_34_17_n_118) | ((mul_34_17_n_6301 & mul_34_17_n_63)
    | (mul_34_17_n_63 & mul_34_17_n_118)));
 assign mul_34_17_n_7600 = (mul_34_17_n_6897 ^ mul_34_17_n_6566);
 assign mul_34_17_n_7795 = ((mul_34_17_n_6128 & mul_34_17_n_6142) | ((mul_34_17_n_6128 & mul_34_17_n_119)
    | (mul_34_17_n_119 & mul_34_17_n_6142)));
 assign mul_34_17_n_7794 = ((mul_34_17_n_6284 & mul_34_17_n_6380) | ((mul_34_17_n_6284 & mul_34_17_n_6285)
    | (mul_34_17_n_6285 & mul_34_17_n_6380)));
 assign mul_34_17_n_7793 = ((mul_34_17_n_6280 & mul_34_17_n_6381) | ((mul_34_17_n_6280 & mul_34_17_n_6281)
    | (mul_34_17_n_6281 & mul_34_17_n_6381)));
 assign mul_34_17_n_7792 = ((mul_34_17_n_6271 & mul_34_17_n_6382) | ((mul_34_17_n_6271 & mul_34_17_n_6273)
    | (mul_34_17_n_6273 & mul_34_17_n_6382)));
 assign mul_34_17_n_7791 = ((mul_34_17_n_6402 & mul_34_17_n_6074) | ((mul_34_17_n_6402 & mul_34_17_n_6682)
    | (mul_34_17_n_6682 & mul_34_17_n_6074)));
 assign mul_34_17_n_7788 = ((mul_34_17_n_6586 & mul_34_17_n_6627) | ((mul_34_17_n_6586 & mul_34_17_n_5710)
    | (mul_34_17_n_5710 & mul_34_17_n_6627)));
 assign mul_34_17_n_7787 = ((mul_34_17_n_6136 & mul_34_17_n_6145) | ((mul_34_17_n_6136 & mul_34_17_n_5116)
    | (mul_34_17_n_5116 & mul_34_17_n_6145)));
 assign mul_34_17_n_7786 = ((mul_34_17_n_6342 & mul_34_17_n_6) | ((mul_34_17_n_6342 & mul_34_17_n_6341)
    | (mul_34_17_n_6341 & mul_34_17_n_6)));
 assign mul_34_17_n_7785 = ((mul_34_17_n_6455 & mul_34_17_n_6511) | ((mul_34_17_n_6455 & mul_34_17_n_6531)
    | (mul_34_17_n_6531 & mul_34_17_n_6511)));
 assign mul_34_17_n_7784 = ((mul_34_17_n_6411 & mul_34_17_n_6424) | ((mul_34_17_n_6411 & mul_34_17_n_5911)
    | (mul_34_17_n_5911 & mul_34_17_n_6424)));
 assign mul_34_17_n_7783 = ((mul_34_17_n_144 & mul_34_17_n_143) | ((mul_34_17_n_144 & mul_34_17_n_5645)
    | (mul_34_17_n_5645 & mul_34_17_n_143)));
 assign mul_34_17_n_7782 = ((mul_34_17_n_6259 & mul_34_17_n_6385) | ((mul_34_17_n_6259 & mul_34_17_n_6254)
    | (mul_34_17_n_6254 & mul_34_17_n_6385)));
 assign mul_34_17_n_7781 = ((mul_34_17_n_17 & mul_34_17_n_12) | ((mul_34_17_n_17 & mul_34_17_n_5122)
    | (mul_34_17_n_5122 & mul_34_17_n_12)));
 assign mul_34_17_n_7779 = ~(mul_34_17_n_6841 ^ mul_34_17_n_5611);
 assign mul_34_17_n_7778 = ((mul_34_17_n_6527 & mul_34_17_n_6626) | ((mul_34_17_n_6527 & mul_34_17_n_6624)
    | (mul_34_17_n_6624 & mul_34_17_n_6626)));
 assign mul_34_17_n_7777 = ((mul_34_17_n_6533 & mul_34_17_n_6640) | ((mul_34_17_n_6533 & mul_34_17_n_6534)
    | (mul_34_17_n_6534 & mul_34_17_n_6640)));
 assign mul_34_17_n_7776 = ((mul_34_17_n_6556 & mul_34_17_n_6668) | ((mul_34_17_n_6556 & mul_34_17_n_6557)
    | (mul_34_17_n_6557 & mul_34_17_n_6668)));
 assign mul_34_17_n_7775 = ((mul_34_17_n_6469 & mul_34_17_n_6512) | ((mul_34_17_n_6469 & mul_34_17_n_6608)
    | (mul_34_17_n_6608 & mul_34_17_n_6512)));
 assign mul_34_17_n_7773 = ~(mul_34_17_n_6912 ^ mul_34_17_n_5512);
 assign mul_34_17_n_7772 = ((mul_34_17_n_6617 & mul_34_17_n_6505) | ((mul_34_17_n_6617 & mul_34_17_n_6480)
    | (mul_34_17_n_6480 & mul_34_17_n_6505)));
 assign mul_34_17_n_7771 = ~(mul_34_17_n_6818 ^ mul_34_17_n_5650);
 assign mul_34_17_n_7770 = ((mul_34_17_n_111 & mul_34_17_n_101) | ((mul_34_17_n_111 & mul_34_17_n_112)
    | (mul_34_17_n_112 & mul_34_17_n_101)));
 assign mul_34_17_n_7769 = ~(mul_34_17_n_6898 ^ mul_34_17_n_19);
 assign mul_34_17_n_7768 = ~(mul_34_17_n_6886 | (mul_34_17_n_6876 | (mul_34_17_n_6118 | mul_34_17_n_4883)));
 assign mul_34_17_n_7767 = ((mul_34_17_n_6584 & mul_34_17_n_6655) | ((mul_34_17_n_6584 & mul_34_17_n_6581)
    | (mul_34_17_n_6581 & mul_34_17_n_6655)));
 assign mul_34_17_n_7766 = ((mul_34_17_n_6306 & mul_34_17_n_6366) | ((mul_34_17_n_6306 & mul_34_17_n_6313)
    | (mul_34_17_n_6313 & mul_34_17_n_6366)));
 assign mul_34_17_n_7765 = ((mul_34_17_n_6219 & mul_34_17_n_6367) | ((mul_34_17_n_6219 & mul_34_17_n_3)
    | (mul_34_17_n_3 & mul_34_17_n_6367)));
 assign mul_34_17_n_7764 = ((mul_34_17_n_6262 & mul_34_17_n_6387) | ((mul_34_17_n_6262 & mul_34_17_n_6261)
    | (mul_34_17_n_6261 & mul_34_17_n_6387)));
 assign mul_34_17_n_7763 = ((mul_34_17_n_6220 & mul_34_17_n_11) | ((mul_34_17_n_6220 & mul_34_17_n_6222)
    | (mul_34_17_n_6222 & mul_34_17_n_11)));
 assign mul_34_17_n_7762 = ((mul_34_17_n_6243 & mul_34_17_n_152) | ((mul_34_17_n_6243 & mul_34_17_n_6240)
    | (mul_34_17_n_6240 & mul_34_17_n_152)));
 assign mul_34_17_n_7761 = ((mul_34_17_n_6298 & mul_34_17_n_5681) | ((mul_34_17_n_6298 & mul_34_17_n_5521)
    | (mul_34_17_n_5521 & mul_34_17_n_5681)));
 assign mul_34_17_n_7760 = ((mul_34_17_n_6585 & mul_34_17_n_58) | ((mul_34_17_n_6585 & mul_34_17_n_5698)
    | (mul_34_17_n_5698 & mul_34_17_n_58)));
 assign mul_34_17_n_7759 = ~((mul_34_17_n_6486 & mul_34_17_n_6573) | (mul_34_17_n_6887 & mul_34_17_n_6517));
 assign mul_34_17_n_7758 = ~(mul_34_17_n_6856 ^ mul_34_17_n_6001);
 assign mul_34_17_n_7757 = ~((mul_34_17_n_6562 & mul_34_17_n_6493) | (mul_34_17_n_6885 & mul_34_17_n_6504));
 assign mul_34_17_n_7756 = ((mul_34_17_n_6129 & mul_34_17_n_6917) | ((mul_34_17_n_6129 & mul_34_17_n_6135)
    | (mul_34_17_n_6135 & mul_34_17_n_6917)));
 assign mul_34_17_n_7754 = ((mul_34_17_n_6546 & mul_34_17_n_190) | ((mul_34_17_n_6546 & mul_34_17_n_6334)
    | (mul_34_17_n_6334 & mul_34_17_n_190)));
 assign mul_34_17_n_7752 = ((mul_34_17_n_6554 & mul_34_17_n_6927) | ((mul_34_17_n_6554 & mul_34_17_n_5921)
    | (mul_34_17_n_5921 & mul_34_17_n_6927)));
 assign mul_34_17_n_7751 = ((mul_34_17_n_6305 & mul_34_17_n_11522) | ((mul_34_17_n_6305 & mul_34_17_n_5)
    | (mul_34_17_n_5 & mul_34_17_n_11522)));
 assign mul_34_17_n_7749 = ((mul_34_17_n_6565 & mul_34_17_n_5884) | ((mul_34_17_n_6565 & mul_34_17_n_5874)
    | (mul_34_17_n_5874 & mul_34_17_n_5884)));
 assign mul_34_17_n_7748 = ((mul_34_17_n_28 & mul_34_17_n_6660) | ((mul_34_17_n_28 & mul_34_17_n_6625)
    | (mul_34_17_n_6625 & mul_34_17_n_6660)));
 assign mul_34_17_n_7747 = ((mul_34_17_n_6248 & mul_34_17_n_6393) | ((mul_34_17_n_6248 & mul_34_17_n_6244)
    | (mul_34_17_n_6244 & mul_34_17_n_6393)));
 assign mul_34_17_n_7746 = ~(mul_34_17_n_6849 ^ mul_34_17_n_5657);
 assign mul_34_17_n_7744 = ((mul_34_17_n_6674 & mul_34_17_n_5798) | ((mul_34_17_n_6674 & mul_34_17_n_6677)
    | (mul_34_17_n_6677 & mul_34_17_n_5798)));
 assign mul_34_17_n_7743 = (mul_34_17_n_6928 ^ mul_34_17_n_5587);
 assign mul_34_17_n_7742 = ((mul_34_17_n_6540 & mul_34_17_n_53) | ((mul_34_17_n_6540 & mul_34_17_n_6535)
    | (mul_34_17_n_6535 & mul_34_17_n_53)));
 assign mul_34_17_n_7741 = ((mul_34_17_n_135 & mul_34_17_n_6684) | ((mul_34_17_n_135 & mul_34_17_n_146)
    | (mul_34_17_n_146 & mul_34_17_n_6684)));
 assign mul_34_17_n_7740 = ((mul_34_17_n_6269 & mul_34_17_n_6202) | ((mul_34_17_n_6269 & mul_34_17_n_6168)
    | (mul_34_17_n_6168 & mul_34_17_n_6202)));
 assign mul_34_17_n_7739 = ((mul_34_17_n_6460 & mul_34_17_n_6516) | ((mul_34_17_n_6460 & mul_34_17_n_6568)
    | (mul_34_17_n_6568 & mul_34_17_n_6516)));
 assign mul_34_17_n_7738 = ~(mul_34_17_n_6847 ^ mul_34_17_n_6029);
 assign mul_34_17_n_7737 = ((mul_34_17_n_6343 & mul_34_17_n_6351) | ((mul_34_17_n_6343 & mul_34_17_n_6265)
    | (mul_34_17_n_6265 & mul_34_17_n_6351)));
 assign mul_34_17_n_7736 = ((mul_34_17_n_6345 & mul_34_17_n_6353) | ((mul_34_17_n_6345 & mul_34_17_n_6346)
    | (mul_34_17_n_6346 & mul_34_17_n_6353)));
 assign mul_34_17_n_7735 = ~(mul_34_17_n_6845 ^ mul_34_17_n_5789);
 assign mul_34_17_n_7734 = ((mul_34_17_n_6412 & mul_34_17_n_6421) | ((mul_34_17_n_6412 & mul_34_17_n_5649)
    | (mul_34_17_n_5649 & mul_34_17_n_6421)));
 assign mul_34_17_n_7733 = ((mul_34_17_n_6547 & mul_34_17_n_6670) | ((mul_34_17_n_6547 & mul_34_17_n_6456)
    | (mul_34_17_n_6456 & mul_34_17_n_6670)));
 assign mul_34_17_n_7732 = ~(mul_34_17_n_6844 ^ mul_34_17_n_5791);
 assign mul_34_17_n_7731 = ((mul_34_17_n_6653 & mul_34_17_n_6506) | ((mul_34_17_n_6653 & mul_34_17_n_6464)
    | (mul_34_17_n_6464 & mul_34_17_n_6506)));
 assign mul_34_17_n_7730 = ~(mul_34_17_n_6843 ^ mul_34_17_n_5624);
 assign mul_34_17_n_7728 = ~(mul_34_17_n_6827 ^ mul_34_17_n_5617);
 assign mul_34_17_n_7727 = ((mul_34_17_n_42 & mul_34_17_n_48) | ((mul_34_17_n_42 & mul_34_17_n_24) |
    (mul_34_17_n_24 & mul_34_17_n_48)));
 assign mul_34_17_n_7726 = ((mul_34_17_n_6536 & mul_34_17_n_6632) | ((mul_34_17_n_6536 & mul_34_17_n_6539)
    | (mul_34_17_n_6539 & mul_34_17_n_6632)));
 assign mul_34_17_n_7725 = ~(mul_34_17_n_6838 ^ mul_34_17_n_6107);
 assign mul_34_17_n_7724 = ~(mul_34_17_n_6837 ^ mul_34_17_n_5792);
 assign mul_34_17_n_7723 = ~(mul_34_17_n_6836 ^ mul_34_17_n_5783);
 assign mul_34_17_n_7722 = ((mul_34_17_n_6320 & mul_34_17_n_6358) | ((mul_34_17_n_6320 & mul_34_17_n_6322)
    | (mul_34_17_n_6322 & mul_34_17_n_6358)));
 assign mul_34_17_n_7720 = ((mul_34_17_n_6544 & mul_34_17_n_107) | ((mul_34_17_n_6544 & mul_34_17_n_6545)
    | (mul_34_17_n_6545 & mul_34_17_n_107)));
 assign mul_34_17_n_7719 = ((mul_34_17_n_6593 & mul_34_17_n_6648) | ((mul_34_17_n_6593 & mul_34_17_n_6591)
    | (mul_34_17_n_6591 & mul_34_17_n_6648)));
 assign mul_34_17_n_7717 = ((mul_34_17_n_6636 & mul_34_17_n_5517) | ((mul_34_17_n_6636 & mul_34_17_n_5509)
    | (mul_34_17_n_5509 & mul_34_17_n_5517)));
 assign mul_34_17_n_7716 = ~(mul_34_17_n_6831 ^ mul_34_17_n_5589);
 assign mul_34_17_n_7715 = ((mul_34_17_n_6467 & mul_34_17_n_6521) | ((mul_34_17_n_6467 & mul_34_17_n_6606)
    | (mul_34_17_n_6606 & mul_34_17_n_6521)));
 assign mul_34_17_n_7714 = ((mul_34_17_n_6471 & mul_34_17_n_2) | ((mul_34_17_n_6471 & mul_34_17_n_6631)
    | (mul_34_17_n_6631 & mul_34_17_n_2)));
 assign mul_34_17_n_7713 = ((mul_34_17_n_6599 & mul_34_17_n_87) | ((mul_34_17_n_6599 & mul_34_17_n_80)
    | (mul_34_17_n_80 & mul_34_17_n_87)));
 assign mul_34_17_n_7712 = ((mul_34_17_n_6329 & mul_34_17_n_150) | ((mul_34_17_n_6329 & mul_34_17_n_6330)
    | (mul_34_17_n_6330 & mul_34_17_n_150)));
 assign mul_34_17_n_7711 = ~(mul_34_17_n_6829 ^ mul_34_17_n_5785);
 assign mul_34_17_n_7710 = ((mul_34_17_n_6472 & mul_34_17_n_6526) | ((mul_34_17_n_6472 & mul_34_17_n_6619)
    | (mul_34_17_n_6619 & mul_34_17_n_6526)));
 assign mul_34_17_n_7708 = ((mul_34_17_n_6594 & mul_34_17_n_82) | ((mul_34_17_n_6594 & mul_34_17_n_6646)
    | (mul_34_17_n_6646 & mul_34_17_n_82)));
 assign mul_34_17_n_7707 = ((mul_34_17_n_6474 & mul_34_17_n_6514) | ((mul_34_17_n_6474 & mul_34_17_n_6623)
    | (mul_34_17_n_6623 & mul_34_17_n_6514)));
 assign mul_34_17_n_7706 = ~(mul_34_17_n_6825 ^ mul_34_17_n_5776);
 assign mul_34_17_n_7705 = ((mul_34_17_n_6478 & mul_34_17_n_6510) | ((mul_34_17_n_6478 & mul_34_17_n_6620)
    | (mul_34_17_n_6620 & mul_34_17_n_6510)));
 assign mul_34_17_n_7704 = ((mul_34_17_n_6294 & mul_34_17_n_6371) | ((mul_34_17_n_6294 & mul_34_17_n_6291)
    | (mul_34_17_n_6291 & mul_34_17_n_6371)));
 assign mul_34_17_n_7703 = ((mul_34_17_n_6489 & mul_34_17_n_6666) | ((mul_34_17_n_6489 & mul_34_17_n_62)
    | (mul_34_17_n_62 & mul_34_17_n_6666)));
 assign mul_34_17_n_7702 = ((mul_34_17_n_6609 & mul_34_17_n_64) | ((mul_34_17_n_6609 & mul_34_17_n_123)
    | (mul_34_17_n_123 & mul_34_17_n_64)));
 assign mul_34_17_n_7701 = ~(mul_34_17_n_6822 ^ mul_34_17_n_133);
 assign mul_34_17_n_7700 = ~(mul_34_17_n_6820 ^ mul_34_17_n_5782);
 assign mul_34_17_n_7699 = ~(mul_34_17_n_6819 ^ mul_34_17_n_6000);
 assign mul_34_17_n_7698 = ~(mul_34_17_n_6850 ^ mul_34_17_n_6023);
 assign mul_34_17_n_7697 = ((mul_34_17_n_6601 & mul_34_17_n_5769) | ((mul_34_17_n_6601 & mul_34_17_n_6602)
    | (mul_34_17_n_6602 & mul_34_17_n_5769)));
 assign mul_34_17_n_7696 = ~(mul_34_17_n_6816 ^ mul_34_17_n_5767);
 assign mul_34_17_n_7695 = ((mul_34_17_n_6588 & mul_34_17_n_6507) | ((mul_34_17_n_6588 & mul_34_17_n_6484)
    | (mul_34_17_n_6484 & mul_34_17_n_6507)));
 assign mul_34_17_n_7694 = ~(mul_34_17_n_6830 ^ mul_34_17_n_5655);
 assign mul_34_17_n_7693 = ((mul_34_17_n_6160 & mul_34_17_n_6628) | ((mul_34_17_n_6160 & mul_34_17_n_6163)
    | (mul_34_17_n_6163 & mul_34_17_n_6628)));
 assign mul_34_17_n_7692 = ((mul_34_17_n_6590 & mul_34_17_n_6922) | ((mul_34_17_n_6590 & mul_34_17_n_6589)
    | (mul_34_17_n_6589 & mul_34_17_n_6922)));
 assign mul_34_17_n_7691 = ((mul_34_17_n_6482 & mul_34_17_n_6523) | ((mul_34_17_n_6482 & mul_34_17_n_6598)
    | (mul_34_17_n_6598 & mul_34_17_n_6523)));
 assign mul_34_17_n_7690 = (mul_34_17_n_6929 ^ mul_34_17_n_6031);
 assign mul_34_17_n_7689 = (mul_34_17_n_6930 ^ mul_34_17_n_6028);
 assign mul_34_17_n_7688 = ((mul_34_17_n_6296 & mul_34_17_n_6398) | ((mul_34_17_n_6296 & mul_34_17_n_6326)
    | (mul_34_17_n_6326 & mul_34_17_n_6398)));
 assign mul_34_17_n_7687 = ((mul_34_17_n_6548 & mul_34_17_n_6671) | ((mul_34_17_n_6548 & mul_34_17_n_6550)
    | (mul_34_17_n_6550 & mul_34_17_n_6671)));
 assign mul_34_17_n_7686 = ~(mul_34_17_n_6846 ^ mul_34_17_n_5697);
 assign mul_34_17_n_7685 = ((mul_34_17_n_38 & mul_34_17_n_6638) | ((mul_34_17_n_38 & mul_34_17_n_41)
    | (mul_34_17_n_41 & mul_34_17_n_6638)));
 assign mul_34_17_n_7684 = ((mul_34_17_n_6537 & mul_34_17_n_6683) | ((mul_34_17_n_6537 & mul_34_17_n_6553)
    | (mul_34_17_n_6553 & mul_34_17_n_6683)));
 assign mul_34_17_n_7682 = ((mul_34_17_n_6325 & mul_34_17_n_6365) | ((mul_34_17_n_6325 & mul_34_17_n_6319)
    | (mul_34_17_n_6319 & mul_34_17_n_6365)));
 assign mul_34_17_n_7680 = ((mul_34_17_n_6338 & mul_34_17_n_6807) | ((mul_34_17_n_6338 & mul_34_17_n_5920)
    | (mul_34_17_n_5920 & mul_34_17_n_6807)));
 assign mul_34_17_n_7679 = ((mul_34_17_n_6347 & mul_34_17_n_6349) | ((mul_34_17_n_6347 & mul_34_17_n_6344)
    | (mul_34_17_n_6344 & mul_34_17_n_6349)));
 assign mul_34_17_n_7678 = ((mul_34_17_n_6415 & mul_34_17_n_6659) | ((mul_34_17_n_6415 & mul_34_17_n_6414)
    | (mul_34_17_n_6414 & mul_34_17_n_6659)));
 assign mul_34_17_n_7677 = ((mul_34_17_n_6237 & mul_34_17_n_5141) | ((mul_34_17_n_6237 & mul_34_17_n_25)
    | (mul_34_17_n_25 & mul_34_17_n_5141)));
 assign mul_34_17_n_7674 = ((mul_34_17_n_6287 & mul_34_17_n_6374) | ((mul_34_17_n_6287 & mul_34_17_n_6289)
    | (mul_34_17_n_6289 & mul_34_17_n_6374)));
 assign mul_34_17_n_7673 = ~(mul_34_17_n_6852 ^ mul_34_17_n_5684);
 assign mul_34_17_n_7671 = ((mul_34_17_n_18 & mul_34_17_n_23) | ((mul_34_17_n_18 & mul_34_17_n_6275)
    | (mul_34_17_n_6275 & mul_34_17_n_23)));
 assign mul_34_17_n_7670 = ~(mul_34_17_n_6824 ^ mul_34_17_n_6105);
 assign mul_34_17_n_7669 = ((mul_34_17_n_6622 & mul_34_17_n_6664) | ((mul_34_17_n_6622 & mul_34_17_n_6621)
    | (mul_34_17_n_6621 & mul_34_17_n_6664)));
 assign mul_34_17_n_7668 = ((mul_34_17_n_6538 & mul_34_17_n_6685) | ((mul_34_17_n_6538 & mul_34_17_n_6541)
    | (mul_34_17_n_6541 & mul_34_17_n_6685)));
 assign mul_34_17_n_7667 = ((mul_34_17_n_6613 & mul_34_17_n_6657) | ((mul_34_17_n_6613 & mul_34_17_n_6019)
    | (mul_34_17_n_6019 & mul_34_17_n_6657)));
 assign mul_34_17_n_7666 = ((mul_34_17_n_117 & mul_34_17_n_66) | ((mul_34_17_n_117 & mul_34_17_n_65)
    | (mul_34_17_n_65 & mul_34_17_n_66)));
 assign mul_34_17_n_7577 = ~mul_34_17_n_7576;
 assign mul_34_17_n_7563 = ~mul_34_17_n_7562;
 assign mul_34_17_n_7558 = ~mul_34_17_n_7557;
 assign mul_34_17_n_7520 = ~mul_34_17_n_7519;
 assign mul_34_17_n_7515 = ~mul_34_17_n_7514;
 assign mul_34_17_n_7505 = ~mul_34_17_n_7504;
 assign mul_34_17_n_7497 = ~mul_34_17_n_7496;
 assign mul_34_17_n_7475 = ~mul_34_17_n_7474;
 assign mul_34_17_n_7472 = ~mul_34_17_n_7471;
 assign mul_34_17_n_7470 = ~mul_34_17_n_158;
 assign mul_34_17_n_7463 = ~mul_34_17_n_7462;
 assign mul_34_17_n_7453 = ~mul_34_17_n_7452;
 assign mul_34_17_n_7449 = ~mul_34_17_n_7448;
 assign mul_34_17_n_7435 = ~mul_34_17_n_7434;
 assign mul_34_17_n_7428 = ~mul_34_17_n_7427;
 assign mul_34_17_n_7422 = ~mul_34_17_n_7421;
 assign mul_34_17_n_7415 = ~mul_34_17_n_7416;
 assign mul_34_17_n_7405 = ~(mul_34_17_n_6795 ^ mul_34_17_n_5516);
 assign mul_34_17_n_7404 = ~(mul_34_17_n_376 | mul_34_17_n_5827);
 assign mul_34_17_n_7403 = ~(mul_34_17_n_6604 ^ mul_34_17_n_6908);
 assign mul_34_17_n_7599 = ~(mul_34_17_n_6744 ^ mul_34_17_n_5763);
 assign mul_34_17_n_7402 = ~(mul_34_17_n_6253 ^ mul_34_17_n_6783);
 assign mul_34_17_n_7598 = ((mul_34_17_n_6152 | mul_34_17_n_5521) & (mul_34_17_n_209 | mul_34_17_n_5681));
 assign mul_34_17_n_7597 = ~(mul_34_17_n_6715 ^ mul_34_17_n_6298);
 assign mul_34_17_n_7401 = (mul_34_17_n_6918 ^ mul_34_17_n_6528);
 assign mul_34_17_n_7400 = (mul_34_17_n_6920 ^ mul_34_17_n_22);
 assign mul_34_17_n_7596 = (mul_34_17_n_6781 ^ mul_34_17_n_27);
 assign mul_34_17_n_7399 = (mul_34_17_n_6532 ^ mul_34_17_n_6777);
 assign mul_34_17_n_7595 = ((mul_34_17_n_6416 & mul_34_17_n_6422) | ((mul_34_17_n_6416 & mul_34_17_n_5654)
    | (mul_34_17_n_5654 & mul_34_17_n_6422)));
 assign mul_34_17_n_7397 = (mul_34_17_n_6786 ^ mul_34_17_n_5968);
 assign mul_34_17_n_7594 = ((mul_34_17_n_6552 & mul_34_17_n_6111) | ((mul_34_17_n_6552 & mul_34_17_n_6618)
    | (mul_34_17_n_6618 & mul_34_17_n_6111)));
 assign mul_34_17_n_7593 = ~(mul_34_17_n_6792 ^ mul_34_17_n_5506);
 assign mul_34_17_n_7592 = ((mul_34_17_n_6312 & mul_34_17_n_5520) | ((mul_34_17_n_6312 & mul_34_17_n_5870)
    | (mul_34_17_n_5870 & mul_34_17_n_5520)));
 assign mul_34_17_n_7591 = ((mul_34_17_n_6221 & mul_34_17_n_6214) | ((mul_34_17_n_6221 & mul_34_17_n_6191)
    | (mul_34_17_n_6191 & mul_34_17_n_6214)));
 assign mul_34_17_n_7590 = ((mul_34_17_n_96 & mul_34_17_n_13) | ((mul_34_17_n_96 & mul_34_17_n_6233)
    | (mul_34_17_n_6233 & mul_34_17_n_13)));
 assign mul_34_17_n_7589 = ~((mul_34_17_n_6934 & ~mul_34_17_n_6368) | (mul_34_17_n_6812 & mul_34_17_n_6368));
 assign mul_34_17_n_7588 = ((mul_34_17_n_6235 & mul_34_17_n_5718) | ((mul_34_17_n_6235 & mul_34_17_n_5140)
    | (mul_34_17_n_5140 & mul_34_17_n_5718)));
 assign mul_34_17_n_7587 = ~(mul_34_17_n_6907 ^ mul_34_17_n_5510);
 assign mul_34_17_n_7586 = ((mul_34_17_n_6161 & mul_34_17_n_6141) | ((mul_34_17_n_6161 & mul_34_17_n_6130)
    | (mul_34_17_n_6130 & mul_34_17_n_6141)));
 assign mul_34_17_n_7585 = ((mul_34_17_n_6165 & mul_34_17_n_6208) | ((mul_34_17_n_6165 & mul_34_17_n_6252)
    | (mul_34_17_n_6252 & mul_34_17_n_6208)));
 assign mul_34_17_n_7584 = ~(mul_34_17_n_6793 ^ mul_34_17_n_6203);
 assign mul_34_17_n_7583 = ~((mul_34_17_n_5886 & (~mul_34_17_n_5505 & ~mul_34_17_n_5119)) | ((mul_34_17_n_5885
    & (mul_34_17_n_5505 & ~mul_34_17_n_5119)) | (mul_34_17_n_6767 & mul_34_17_n_5119)));
 assign mul_34_17_n_7582 = ((mul_34_17_n_6189 & mul_34_17_n_6205) | ((mul_34_17_n_6189 & mul_34_17_n_6266)
    | (mul_34_17_n_6266 & mul_34_17_n_6205)));
 assign mul_34_17_n_7581 = ~(mul_34_17_n_6701 ^ mul_34_17_n_5575);
 assign mul_34_17_n_7580 = ~(mul_34_17_n_6707 ^ mul_34_17_n_6010);
 assign mul_34_17_n_7579 = ~(mul_34_17_n_6711 ^ mul_34_17_n_5584);
 assign mul_34_17_n_7576 = ((mul_34_17_n_6654 & mul_34_17_n_91) | ((mul_34_17_n_6654 & mul_34_17_n_81)
    | (mul_34_17_n_81 & mul_34_17_n_91)));
 assign mul_34_17_n_7573 = ~((mul_34_17_n_2810 & (~mul_34_17_n_5431 & ~mul_34_17_n_6848)) | ((mul_34_17_n_2809
    & (mul_34_17_n_5431 & ~mul_34_17_n_6848)) | (mul_34_17_n_6681 & mul_34_17_n_6848)));
 assign mul_34_17_n_7572 = ((mul_34_17_n_6871 & mul_34_17_n_6401) | (mul_34_17_n_6883 & mul_34_17_n_6449));
 assign mul_34_17_n_7570 = ~(mul_34_17_n_6795 ^ mul_34_17_n_5515);
 assign mul_34_17_n_7568 = ((mul_34_17_n_6495 & mul_34_17_n_6509) | ((mul_34_17_n_6495 & mul_34_17_n_6542)
    | (mul_34_17_n_6542 & mul_34_17_n_6509)));
 assign mul_34_17_n_7567 = ((mul_34_17_n_6167 & mul_34_17_n_6196) | ((mul_34_17_n_6167 & mul_34_17_n_6328)
    | (mul_34_17_n_6328 & mul_34_17_n_6196)));
 assign mul_34_17_n_7566 = ((mul_34_17_n_6610 & mul_34_17_n_6629) | ((mul_34_17_n_6610 & mul_34_17_n_6614)
    | (mul_34_17_n_6614 & mul_34_17_n_6629)));
 assign mul_34_17_n_7565 = ~(mul_34_17_n_6692 ^ mul_34_17_n_5578);
 assign mul_34_17_n_7564 = ((mul_34_17_n_6355 & mul_34_17_n_6195) | ((mul_34_17_n_6355 & mul_34_17_n_6190)
    | (mul_34_17_n_6190 & mul_34_17_n_6195)));
 assign mul_34_17_n_7562 = ~(mul_34_17_n_6796 ^ mul_34_17_n_5875);
 assign mul_34_17_n_7561 = ~(mul_34_17_n_6733 ^ mul_34_17_n_5673);
 assign mul_34_17_n_7560 = ((mul_34_17_n_6126 & mul_34_17_n_6143) | ((mul_34_17_n_6126 & mul_34_17_n_5706)
    | (mul_34_17_n_5706 & mul_34_17_n_6143)));
 assign mul_34_17_n_7559 = ((mul_34_17_n_6483 & mul_34_17_n_6525) | ((mul_34_17_n_6483 & mul_34_17_n_6644)
    | (mul_34_17_n_6644 & mul_34_17_n_6525)));
 assign mul_34_17_n_7557 = ~(mul_34_17_n_6788 ^ mul_34_17_n_6216);
 assign mul_34_17_n_7556 = ((mul_34_17_n_6156 & mul_34_17_n_6801) | ((mul_34_17_n_6156 & mul_34_17_n_6174)
    | (mul_34_17_n_6174 & mul_34_17_n_6801)));
 assign mul_34_17_n_7555 = ((mul_34_17_n_26 & mul_34_17_n_6369) | ((mul_34_17_n_26 & mul_34_17_n_6286)
    | (mul_34_17_n_6286 & mul_34_17_n_6369)));
 assign mul_34_17_n_7554 = ((mul_34_17_n_6175 & mul_34_17_n_6139) | ((mul_34_17_n_6175 & mul_34_17_n_6125)
    | (mul_34_17_n_6125 & mul_34_17_n_6139)));
 assign mul_34_17_n_7553 = ((mul_34_17_n_55 & mul_34_17_n_39) | ((mul_34_17_n_55 & mul_34_17_n_40) |
    (mul_34_17_n_40 & mul_34_17_n_39)));
 assign mul_34_17_n_7552 = ((mul_34_17_n_6363 & mul_34_17_n_6211) | ((mul_34_17_n_6363 & mul_34_17_n_6159)
    | (mul_34_17_n_6159 & mul_34_17_n_6211)));
 assign mul_34_17_n_7551 = ((mul_34_17_n_6227 & mul_34_17_n_6375) | ((mul_34_17_n_6227 & mul_34_17_n_5630)
    | (mul_34_17_n_5630 & mul_34_17_n_6375)));
 assign mul_34_17_n_7550 = ~(mul_34_17_n_6743 ^ mul_34_17_n_5739);
 assign mul_34_17_n_7549 = ~(mul_34_17_n_6747 ^ mul_34_17_n_5946);
 assign mul_34_17_n_7548 = ~(mul_34_17_n_6754 ^ mul_34_17_n_5958);
 assign mul_34_17_n_7547 = ((mul_34_17_n_6170 & mul_34_17_n_6212) | ((mul_34_17_n_6170 & mul_34_17_n_6230)
    | (mul_34_17_n_6230 & mul_34_17_n_6212)));
 assign mul_34_17_n_7546 = ((mul_34_17_n_6302 & mul_34_17_n_6199) | ((mul_34_17_n_6302 & mul_34_17_n_6303)
    | (mul_34_17_n_6303 & mul_34_17_n_6199)));
 assign mul_34_17_n_7545 = ~(mul_34_17_n_6746 ^ mul_34_17_n_5917);
 assign mul_34_17_n_7544 = ~(mul_34_17_n_6745 ^ mul_34_17_n_5712);
 assign mul_34_17_n_7542 = ~(mul_34_17_n_6758 ^ mul_34_17_n_6102);
 assign mul_34_17_n_7541 = ((mul_34_17_n_6226 & mul_34_17_n_6923) | ((mul_34_17_n_6226 & mul_34_17_n_6224)
    | (mul_34_17_n_6224 & mul_34_17_n_6923)));
 assign mul_34_17_n_7540 = ((mul_34_17_n_6278 & mul_34_17_n_6630) | ((mul_34_17_n_6278 & mul_34_17_n_5988)
    | (mul_34_17_n_5988 & mul_34_17_n_6630)));
 assign mul_34_17_n_7539 = ~(mul_34_17_n_5966 ^ mul_34_17_n_6757);
 assign mul_34_17_n_7538 = ((mul_34_17_n_6564 & mul_34_17_n_6919) | ((mul_34_17_n_6564 & mul_34_17_n_115)
    | (mul_34_17_n_115 & mul_34_17_n_6919)));
 assign mul_34_17_n_7537 = ~(mul_34_17_n_6741 ^ mul_34_17_n_5120);
 assign mul_34_17_n_7536 = ((mul_34_17_n_6529 & mul_34_17_n_6663) | ((mul_34_17_n_6529 & mul_34_17_n_5669)
    | (mul_34_17_n_5669 & mul_34_17_n_6663)));
 assign mul_34_17_n_7535 = ~(mul_34_17_n_6730 ^ mul_34_17_n_99);
 assign mul_34_17_n_7534 = ~(mul_34_17_n_6739 ^ mul_34_17_n_6101);
 assign mul_34_17_n_7533 = ~(mul_34_17_n_6737 ^ mul_34_17_n_6050);
 assign mul_34_17_n_7532 = ((mul_34_17_n_6642 & mul_34_17_n_6501) | ((mul_34_17_n_6642 & mul_34_17_n_6481)
    | (mul_34_17_n_6481 & mul_34_17_n_6501)));
 assign mul_34_17_n_7531 = ~(mul_34_17_n_6693 ^ mul_34_17_n_5779);
 assign mul_34_17_n_7530 = ((mul_34_17_n_6419 & mul_34_17_n_6420) | ((mul_34_17_n_6419 & mul_34_17_n_6635)
    | (mul_34_17_n_6635 & mul_34_17_n_6420)));
 assign mul_34_17_n_7529 = ~(mul_34_17_n_6734 ^ mul_34_17_n_5546);
 assign mul_34_17_n_7528 = ~(mul_34_17_n_6810 ^ mul_34_17_n_5582);
 assign mul_34_17_n_7527 = ((mul_34_17_n_6354 & mul_34_17_n_6197) | ((mul_34_17_n_6354 & mul_34_17_n_6169)
    | (mul_34_17_n_6169 & mul_34_17_n_6197)));
 assign mul_34_17_n_7526 = ((mul_34_17_n_6336 & mul_34_17_n_6360) | ((mul_34_17_n_6336 & mul_34_17_n_6186)
    | (mul_34_17_n_6186 & mul_34_17_n_6360)));
 assign mul_34_17_n_7525 = ~(mul_34_17_n_6811 ^ mul_34_17_n_5574);
 assign mul_34_17_n_7524 = ((mul_34_17_n_14 & mul_34_17_n_51) | ((mul_34_17_n_14 & mul_34_17_n_45) |
    (mul_34_17_n_45 & mul_34_17_n_51)));
 assign mul_34_17_n_7523 = ~(mul_34_17_n_6760 ^ mul_34_17_n_5967);
 assign mul_34_17_n_7522 = ~(mul_34_17_n_6729 ^ mul_34_17_n_89);
 assign mul_34_17_n_7521 = ((mul_34_17_n_6576 & mul_34_17_n_6524) | ((mul_34_17_n_6576 & mul_34_17_n_5412)
    | (mul_34_17_n_5412 & mul_34_17_n_6524)));
 assign mul_34_17_n_7519 = ~(mul_34_17_n_6728 ^ mul_34_17_n_6067);
 assign mul_34_17_n_7518 = ((mul_34_17_n_6324 & mul_34_17_n_6357) | ((mul_34_17_n_6324 & mul_34_17_n_73)
    | (mul_34_17_n_73 & mul_34_17_n_6357)));
 assign mul_34_17_n_7517 = ~(mul_34_17_n_6727 ^ mul_34_17_n_5690);
 assign mul_34_17_n_7516 = ~(mul_34_17_n_6698 ^ mul_34_17_n_5732);
 assign mul_34_17_n_7514 = ((mul_34_17_n_6282 & mul_34_17_n_97) | ((mul_34_17_n_6282 & mul_34_17_n_79)
    | (mul_34_17_n_79 & mul_34_17_n_97)));
 assign mul_34_17_n_7513 = ~(mul_34_17_n_6763 ^ mul_34_17_n_5970);
 assign mul_34_17_n_7512 = ((mul_34_17_n_6348 & mul_34_17_n_6384) | ((mul_34_17_n_6348 & mul_34_17_n_6162)
    | (mul_34_17_n_6162 & mul_34_17_n_6384)));
 assign mul_34_17_n_7511 = ~(mul_34_17_n_6109 ^ (mul_34_17_n_5992 ^ (mul_34_17_n_4829 ^ mul_34_17_n_4828)));
 assign mul_34_17_n_7509 = ((mul_34_17_n_6332 & mul_34_17_n_6192) | ((mul_34_17_n_6332 & mul_34_17_n_6153)
    | (mul_34_17_n_6153 & mul_34_17_n_6192)));
 assign mul_34_17_n_7508 = ((mul_34_17_n_88 & mul_34_17_n_6397) | ((mul_34_17_n_88 & mul_34_17_n_98)
    | (mul_34_17_n_98 & mul_34_17_n_6397)));
 assign mul_34_17_n_7507 = ~(mul_34_17_n_6718 ^ mul_34_17_n_5533);
 assign mul_34_17_n_7506 = ~(mul_34_17_n_6722 ^ mul_34_17_n_5680);
 assign mul_34_17_n_7396 = ~(mul_34_17_n_6809 ^ mul_34_17_n_5620);
 assign mul_34_17_n_7395 = (mul_34_17_n_6806 ^ mul_34_17_n_5586);
 assign mul_34_17_n_7504 = ((mul_34_17_n_6132 & mul_34_17_n_6508) | ((mul_34_17_n_6132 & mul_34_17_n_6133)
    | (mul_34_17_n_6133 & mul_34_17_n_6508)));
 assign mul_34_17_n_7503 = ~(mul_34_17_n_6713 ^ mul_34_17_n_85);
 assign mul_34_17_n_7501 = ((mul_34_17_n_92 & mul_34_17_n_6201) | ((mul_34_17_n_92 & mul_34_17_n_52)
    | (mul_34_17_n_52 & mul_34_17_n_6201)));
 assign mul_34_17_n_7500 = ~(mul_34_17_n_6720 ^ mul_34_17_n_5579);
 assign mul_34_17_n_7499 = ((mul_34_17_n_102 & mul_34_17_n_6425) | ((mul_34_17_n_102 & mul_34_17_n_6131)
    | (mul_34_17_n_6131 & mul_34_17_n_6425)));
 assign mul_34_17_n_7498 = ~(mul_34_17_n_6710 ^ mul_34_17_n_5608);
 assign mul_34_17_n_7496 = ~(mul_34_17_n_6709 ^ mul_34_17_n_5682);
 assign mul_34_17_n_7495 = ((mul_34_17_n_6290 & mul_34_17_n_6373) | ((mul_34_17_n_6290 & mul_34_17_n_6172)
    | (mul_34_17_n_6172 & mul_34_17_n_6373)));
 assign mul_34_17_n_7494 = ((mul_34_17_n_6579 & mul_34_17_n_95) | ((mul_34_17_n_6579 & mul_34_17_n_20)
    | (mul_34_17_n_20 & mul_34_17_n_95)));
 assign mul_34_17_n_7493 = ~(mul_34_17_n_6842 ^ mul_34_17_n_5518);
 assign mul_34_17_n_7492 = ~(mul_34_17_n_6860 ^ mul_34_17_n_5665);
 assign mul_34_17_n_7491 = ~(mul_34_17_n_6705 ^ mul_34_17_n_6081);
 assign mul_34_17_n_7490 = ((mul_34_17_n_19 & mul_34_17_n_5764) | ((mul_34_17_n_19 & mul_34_17_n_5689)
    | (mul_34_17_n_5689 & mul_34_17_n_5764)));
 assign mul_34_17_n_7489 = ~(mul_34_17_n_6704 ^ mul_34_17_n_5588);
 assign mul_34_17_n_7488 = ~(mul_34_17_n_6703 ^ mul_34_17_n_5685);
 assign mul_34_17_n_7487 = ((mul_34_17_n_6283 & mul_34_17_n_6379) | ((mul_34_17_n_6283 & mul_34_17_n_5568)
    | (mul_34_17_n_5568 & mul_34_17_n_6379)));
 assign mul_34_17_n_7486 = ~(mul_34_17_n_6702 ^ mul_34_17_n_5570);
 assign mul_34_17_n_7484 = ~(mul_34_17_n_6700 ^ mul_34_17_n_5563);
 assign mul_34_17_n_7483 = ~(mul_34_17_n_6699 ^ mul_34_17_n_5758);
 assign mul_34_17_n_7482 = ((mul_34_17_n_6267 & mul_34_17_n_6204) | ((mul_34_17_n_6267 & mul_34_17_n_6164)
    | (mul_34_17_n_6164 & mul_34_17_n_6204)));
 assign mul_34_17_n_7481 = ((mul_34_17_n_6543 & mul_34_17_n_6520) | ((mul_34_17_n_6543 & mul_34_17_n_6607)
    | (mul_34_17_n_6607 & mul_34_17_n_6520)));
 assign mul_34_17_n_7480 = ((mul_34_17_n_6166 & mul_34_17_n_6209) | ((mul_34_17_n_6166 & mul_34_17_n_6390)
    | (mul_34_17_n_6390 & mul_34_17_n_6209)));
 assign mul_34_17_n_7479 = ((mul_34_17_n_6256 & mul_34_17_n_6206) | ((mul_34_17_n_6256 & mul_34_17_n_6181)
    | (mul_34_17_n_6181 & mul_34_17_n_6206)));
 assign mul_34_17_n_7478 = ~(mul_34_17_n_6697 ^ mul_34_17_n_6034);
 assign mul_34_17_n_7476 = ((mul_34_17_n_6413 & mul_34_17_n_6426) | ((mul_34_17_n_6413 & mul_34_17_n_6003)
    | (mul_34_17_n_6003 & mul_34_17_n_6426)));
 assign mul_34_17_n_7474 = ~(mul_34_17_n_6695 ^ mul_34_17_n_5111);
 assign mul_34_17_n_7473 = ~(mul_34_17_n_6696 ^ mul_34_17_n_5778);
 assign mul_34_17_n_7471 = ((mul_34_17_n_6225 & mul_34_17_n_6641) | ((mul_34_17_n_6225 & mul_34_17_n_10)
    | (mul_34_17_n_10 & mul_34_17_n_6641)));
 assign mul_34_17_n_7394 = (mul_34_17_n_6803 ^ mul_34_17_n_5552);
 assign mul_34_17_n_7469 = ~(mul_34_17_n_6753 ^ mul_34_17_n_5648);
 assign mul_34_17_n_7468 = ~(mul_34_17_n_6690 ^ mul_34_17_n_5544);
 assign mul_34_17_n_7467 = ((mul_34_17_n_6465 & mul_34_17_n_6639) | ((mul_34_17_n_6465 & mul_34_17_n_6600)
    | (mul_34_17_n_6600 & mul_34_17_n_6639)));
 assign mul_34_17_n_7466 = ~(mul_34_17_n_6712 ^ mul_34_17_n_5564);
 assign mul_34_17_n_7465 = ~(mul_34_17_n_6717 ^ mul_34_17_n_5535);
 assign mul_34_17_n_7393 = ~(mul_34_17_n_6805 ^ mul_34_17_n_5538);
 assign mul_34_17_n_7464 = ((mul_34_17_n_6127 & mul_34_17_n_6144) | ((mul_34_17_n_6127 & mul_34_17_n_5529)
    | (mul_34_17_n_5529 & mul_34_17_n_6144)));
 assign mul_34_17_n_7462 = ((mul_34_17_n_15 & mul_34_17_n_16) | ((mul_34_17_n_15 & mul_34_17_n_5677)
    | (mul_34_17_n_5677 & mul_34_17_n_16)));
 assign mul_34_17_n_7461 = ((mul_34_17_n_6316 & mul_34_17_n_69) | ((mul_34_17_n_6316 & mul_34_17_n_5871)
    | (mul_34_17_n_5871 & mul_34_17_n_69)));
 assign mul_34_17_n_7460 = ((mul_34_17_n_6574 & mul_34_17_n_93) | ((mul_34_17_n_6574 & mul_34_17_n_5947)
    | (mul_34_17_n_5947 & mul_34_17_n_93)));
 assign mul_34_17_n_7459 = ((mul_34_17_n_6183 & mul_34_17_n_6406) | ((mul_34_17_n_6183 & mul_34_17_n_6178)
    | (mul_34_17_n_6178 & mul_34_17_n_6406)));
 assign mul_34_17_n_7458 = ~(mul_34_17_n_6723 ^ mul_34_17_n_5597);
 assign mul_34_17_n_7457 = ((mul_34_17_n_6229 & mul_34_17_n_6370) | ((mul_34_17_n_6229 & mul_34_17_n_6176)
    | (mul_34_17_n_6176 & mul_34_17_n_6370)));
 assign mul_34_17_n_7456 = ~(mul_34_17_n_6749 ^ mul_34_17_n_5522);
 assign mul_34_17_n_7455 = ~(mul_34_17_n_6750 ^ mul_34_17_n_5632);
 assign mul_34_17_n_7454 = ~(mul_34_17_n_6751 ^ mul_34_17_n_5803);
 assign mul_34_17_n_7452 = ((mul_34_17_n_31 & mul_34_17_n_29) | ((mul_34_17_n_31 & mul_34_17_n_30) |
    (mul_34_17_n_30 & mul_34_17_n_29)));
 assign mul_34_17_n_7392 = (mul_34_17_n_6932 ^ mul_34_17_n_6033);
 assign mul_34_17_n_7451 = ((mul_34_17_n_6255 & mul_34_17_n_5802) | ((mul_34_17_n_6255 & mul_34_17_n_6250)
    | (mul_34_17_n_6250 & mul_34_17_n_5802)));
 assign mul_34_17_n_7450 = ~(mul_34_17_n_6756 ^ mul_34_17_n_5596);
 assign mul_34_17_n_7448 = ((mul_34_17_n_6182 & mul_34_17_n_6218) | ((mul_34_17_n_6182 & mul_34_17_n_6223)
    | (mul_34_17_n_6223 & mul_34_17_n_6218)));
 assign mul_34_17_n_7447 = ~(mul_34_17_n_6759 ^ mul_34_17_n_5561);
 assign mul_34_17_n_7391 = ~(mul_34_17_n_6925 ^ mul_34_17_n_6071);
 assign mul_34_17_n_7446 = ~(mul_34_17_n_6764 ^ mul_34_17_n_5772);
 assign mul_34_17_n_7445 = ((mul_34_17_n_6395 & mul_34_17_n_6667) | ((mul_34_17_n_6395 & mul_34_17_n_6270)
    | (mul_34_17_n_6270 & mul_34_17_n_6667)));
 assign mul_34_17_n_7444 = ~(mul_34_17_n_6859 ^ mul_34_17_n_5896);
 assign mul_34_17_n_7443 = ~(mul_34_17_n_6823 ^ mul_34_17_n_5687);
 assign mul_34_17_n_7442 = ((mul_34_17_n_6466 & mul_34_17_n_121) | ((mul_34_17_n_6466 & mul_34_17_n_120)
    | (mul_34_17_n_120 & mul_34_17_n_121)));
 assign mul_34_17_n_7441 = ~(mul_34_17_n_6706 ^ mul_34_17_n_5695);
 assign mul_34_17_n_7440 = ~(mul_34_17_n_6731 ^ mul_34_17_n_5647);
 assign mul_34_17_n_7439 = ((mul_34_17_n_6577 & mul_34_17_n_6499) | ((mul_34_17_n_6577 & mul_34_17_n_6488)
    | (mul_34_17_n_6488 & mul_34_17_n_6499)));
 assign mul_34_17_n_7438 = ~(mul_34_17_n_6821 ^ mul_34_17_n_5757);
 assign mul_34_17_n_7437 = ((mul_34_17_n_6249 & mul_34_17_n_6391) | ((mul_34_17_n_6249 & mul_34_17_n_5118)
    | (mul_34_17_n_5118 & mul_34_17_n_6391)));
 assign mul_34_17_n_7436 = ((mul_34_17_n_6245 & mul_34_17_n_6210) | ((mul_34_17_n_6245 & mul_34_17_n_6154)
    | (mul_34_17_n_6154 & mul_34_17_n_6210)));
 assign mul_34_17_n_7434 = ~(mul_34_17_n_6719 ^ mul_34_17_n_5640);
 assign mul_34_17_n_7433 = ~(mul_34_17_n_6736 ^ mul_34_17_n_5603);
 assign mul_34_17_n_7431 = ((mul_34_17_n_6297 & mul_34_17_n_6198) | ((mul_34_17_n_6297 & mul_34_17_n_5410)
    | (mul_34_17_n_5410 & mul_34_17_n_6198)));
 assign mul_34_17_n_7430 = ((mul_34_17_n_6479 & mul_34_17_n_6518) | ((mul_34_17_n_6479 & mul_34_17_n_6315)
    | (mul_34_17_n_6315 & mul_34_17_n_6518)));
 assign mul_34_17_n_7429 = ((mul_34_17_n_6311 & mul_34_17_n_6215) | ((mul_34_17_n_6311 & mul_34_17_n_6158)
    | (mul_34_17_n_6158 & mul_34_17_n_6215)));
 assign mul_34_17_n_7427 = ((mul_34_17_n_6228 & mul_34_17_n_6399) | ((mul_34_17_n_6228 & mul_34_17_n_5532)
    | (mul_34_17_n_5532 & mul_34_17_n_6399)));
 assign mul_34_17_n_7425 = ~(mul_34_17_n_6735 ^ mul_34_17_n_5602);
 assign mul_34_17_n_7424 = ~(mul_34_17_n_6861 ^ mul_34_17_n_6093);
 assign mul_34_17_n_7423 = ((mul_34_17_n_6246 & mul_34_17_n_6394) | ((mul_34_17_n_6246 & mul_34_17_n_6247)
    | (mul_34_17_n_6247 & mul_34_17_n_6394)));
 assign mul_34_17_n_7421 = ((mul_34_17_n_6317 & mul_34_17_n_6213) | ((mul_34_17_n_6317 & mul_34_17_n_6179)
    | (mul_34_17_n_6179 & mul_34_17_n_6213)));
 assign mul_34_17_n_7420 = ~(mul_34_17_n_6726 ^ mul_34_17_n_5664);
 assign mul_34_17_n_7418 = ~(mul_34_17_n_6738 ^ mul_34_17_n_5900);
 assign mul_34_17_n_7416 = ~(mul_34_17_n_6708 ^ mul_34_17_n_5678);
 assign mul_34_17_n_7414 = ((mul_34_17_n_6452 & mul_34_17_n_6500) | ((mul_34_17_n_6452 & mul_34_17_n_6530)
    | (mul_34_17_n_6530 & mul_34_17_n_6500)));
 assign mul_34_17_n_7413 = ~(mul_34_17_n_6725 ^ mul_34_17_n_5539);
 assign mul_34_17_n_7412 = (mul_34_17_n_6804 ^ mul_34_17_n_5906);
 assign mul_34_17_n_7411 = ~(mul_34_17_n_6721 ^ mul_34_17_n_5731);
 assign mul_34_17_n_7410 = ~(mul_34_17_n_6732 ^ mul_34_17_n_5963);
 assign mul_34_17_n_7408 = ((mul_34_17_n_6335 & mul_34_17_n_6194) | ((mul_34_17_n_6335 & mul_34_17_n_6333)
    | (mul_34_17_n_6333 & mul_34_17_n_6194)));
 assign mul_34_17_n_7407 = ~(mul_34_17_n_6740 ^ mul_34_17_n_5580);
 assign mul_34_17_n_7390 = ~mul_34_17_n_7258;
 assign mul_34_17_n_7389 = ~mul_34_17_n_7251;
 assign mul_34_17_n_7369 = ~mul_34_17_n_7368;
 assign mul_34_17_n_7366 = ~mul_34_17_n_7365;
 assign mul_34_17_n_7357 = ~mul_34_17_n_7356;
 assign mul_34_17_n_7349 = ~mul_34_17_n_7350;
 assign mul_34_17_n_7348 = ~mul_34_17_n_7347;
 assign mul_34_17_n_7329 = ~mul_34_17_n_7328;
 assign mul_34_17_n_7326 = ~mul_34_17_n_7325;
 assign mul_34_17_n_7319 = ~mul_34_17_n_7318;
 assign mul_34_17_n_7316 = ~mul_34_17_n_7315;
 assign mul_34_17_n_7300 = ~mul_34_17_n_7299;
 assign mul_34_17_n_7294 = ~mul_34_17_n_7293;
 assign mul_34_17_n_7289 = ~mul_34_17_n_7290;
 assign mul_34_17_n_7288 = (mul_34_17_n_6499 ^ mul_34_17_n_6488);
 assign mul_34_17_n_7287 = ~(mul_34_17_n_6781 & mul_34_17_n_6299);
 assign mul_34_17_n_7286 = ~(mul_34_17_n_6782 & mul_34_17_n_27);
 assign mul_34_17_n_7285 = ~(mul_34_17_n_6867 | mul_34_17_n_5816);
 assign mul_34_17_n_7284 = (mul_34_17_n_6537 ^ mul_34_17_n_6553);
 assign mul_34_17_n_7283 = ~(mul_34_17_n_389 | mul_34_17_n_5860);
 assign mul_34_17_n_7282 = (mul_34_17_n_6527 ^ mul_34_17_n_6624);
 assign mul_34_17_n_7281 = ~(mul_34_17_n_6864 | mul_34_17_n_5857);
 assign mul_34_17_n_7280 = ~(mul_34_17_n_6329 ^ mul_34_17_n_6330);
 assign mul_34_17_n_7278 = ~(mul_34_17_n_6898 & mul_34_17_n_19);
 assign mul_34_17_n_7277 = ~(mul_34_17_n_6898 | mul_34_17_n_19);
 assign mul_34_17_n_7276 = ~(mul_34_17_n_6910 & mul_34_17_n_5514);
 assign mul_34_17_n_7274 = ~(mul_34_17_n_6408 ^ mul_34_17_n_6687);
 assign mul_34_17_n_7273 = (mul_34_17_n_6544 ^ mul_34_17_n_6545);
 assign mul_34_17_n_7268 = ~(mul_34_17_n_6870 & mul_34_17_n_5850);
 assign mul_34_17_n_7267 = ~(mul_34_17_n_6554 ^ mul_34_17_n_5921);
 assign mul_34_17_n_7266 = ~(mul_34_17_n_6537 ^ mul_34_17_n_6553);
 assign mul_34_17_n_7265 = (mul_34_17_n_6622 ^ mul_34_17_n_6621);
 assign mul_34_17_n_7263 = ~(mul_34_17_n_6791 | mul_34_17_n_5507);
 assign mul_34_17_n_7261 = ~(mul_34_17_n_6788 & mul_34_17_n_6217);
 assign mul_34_17_n_7260 = ~(mul_34_17_n_6788 | mul_34_17_n_6217);
 assign mul_34_17_n_7259 = (mul_34_17_n_6248 ^ mul_34_17_n_6244);
 assign mul_34_17_n_7258 = ~(mul_34_17_n_6792 | mul_34_17_n_5506);
 assign mul_34_17_n_7256 = ~(mul_34_17_n_6343 ^ mul_34_17_n_6265);
 assign mul_34_17_n_7255 = ~(mul_34_17_n_6345 ^ mul_34_17_n_6346);
 assign mul_34_17_n_7253 = (mul_34_17_n_5464 ^ mul_34_17_n_6403);
 assign mul_34_17_n_7252 = ~(mul_34_17_n_6813 & mul_34_17_n_6368);
 assign mul_34_17_n_7251 = ~(mul_34_17_n_6934 | mul_34_17_n_6368);
 assign mul_34_17_n_7250 = ~(mul_34_17_n_6546 ^ mul_34_17_n_6334);
 assign mul_34_17_n_7249 = (mul_34_17_n_6262 ^ mul_34_17_n_6261);
 assign mul_34_17_n_7248 = ~(mul_34_17_n_6793 & mul_34_17_n_6203);
 assign mul_34_17_n_7247 = ~(mul_34_17_n_6793 | mul_34_17_n_6203);
 assign mul_34_17_n_7246 = ~(mul_34_17_n_6183 ^ mul_34_17_n_6178);
 assign mul_34_17_n_7245 = (mul_34_17_n_6220 ^ mul_34_17_n_6222);
 assign mul_34_17_n_7244 = ~(mul_34_17_n_5921 ^ mul_34_17_n_6554);
 assign mul_34_17_n_7242 = ~(mul_34_17_n_6347 ^ mul_34_17_n_6344);
 assign mul_34_17_n_7240 = ~(mul_34_17_n_6195 ^ mul_34_17_n_6190);
 assign mul_34_17_n_7238 = ((mul_34_17_n_5822 & mul_34_17_n_5823) | (mul_34_17_n_6445 & mul_34_17_n_5821));
 assign mul_34_17_n_7237 = ~(mul_34_17_n_5169 ^ (mul_34_17_n_4619 ^ (mul_34_17_n_5453 ^ mul_34_17_n_4620)));
 assign mul_34_17_n_7233 = (mul_34_17_n_6509 ^ mul_34_17_n_6495);
 assign mul_34_17_n_7230 = ~(mul_34_17_n_5455 ^ (mul_34_17_n_4018 ^ (mul_34_17_n_5456 ^ mul_34_17_n_4582)));
 assign mul_34_17_n_7220 = ~(mul_34_17_n_6524 ^ mul_34_17_n_5413);
 assign mul_34_17_n_7219 = ((mul_34_17_n_5820 & mul_34_17_n_5818) | (mul_34_17_n_6431 & mul_34_17_n_5696));
 assign mul_34_17_n_7218 = ~(mul_34_17_n_6482 ^ mul_34_17_n_6523);
 assign mul_34_17_n_7217 = ~(mul_34_17_n_5462 ^ (mul_34_17_n_3591 ^ (mul_34_17_n_5461 ^ mul_34_17_n_4676)));
 assign mul_34_17_n_7216 = ((mul_34_17_n_5826 & mul_34_17_n_5825) | (mul_34_17_n_6433 & mul_34_17_n_5824));
 assign mul_34_17_n_7210 = ~(mul_34_17_n_5481 ^ (mul_34_17_n_2837 ^ (mul_34_17_n_5480 ^ mul_34_17_n_4789)));
 assign mul_34_17_n_7209 = ~(mul_34_17_n_6461 ^ mul_34_17_n_6502);
 assign mul_34_17_n_7208 = ~(mul_34_17_n_5175 ^ (mul_34_17_n_3883 ^ (mul_34_17_n_5170 ^ mul_34_17_n_3100)));
 assign mul_34_17_n_7207 = ~(mul_34_17_n_5467 ^ (mul_34_17_n_4714 ^ (mul_34_17_n_5466 ^ mul_34_17_n_3860)));
 assign mul_34_17_n_7205 = ((mul_34_17_n_5872 & mul_34_17_n_390) | ((mul_34_17_n_5872 & mul_34_17_n_3979)
    | (mul_34_17_n_3979 & mul_34_17_n_390)));
 assign mul_34_17_n_7199 = ~(mul_34_17_n_5185 ^ (mul_34_17_n_3890 ^ (mul_34_17_n_5186 ^ mul_34_17_n_3892)));
 assign mul_34_17_n_7198 = ~(mul_34_17_n_6595 ^ mul_34_17_n_5427);
 assign mul_34_17_n_7195 = ~(mul_34_17_n_6511 ^ mul_34_17_n_145);
 assign mul_34_17_n_7194 = ~(mul_34_17_n_5484 ^ (mul_34_17_n_4791 ^ (mul_34_17_n_5483 ^ mul_34_17_n_4788)));
 assign mul_34_17_n_7193 = (mul_34_17_n_6460 ^ mul_34_17_n_6516);
 assign mul_34_17_n_7191 = ~(mul_34_17_n_6464 ^ mul_34_17_n_6506);
 assign mul_34_17_n_7190 = ~(mul_34_17_n_5479 ^ (mul_34_17_n_3691 ^ (mul_34_17_n_5477 ^ mul_34_17_n_4775)));
 assign mul_34_17_n_7189 = ~(mul_34_17_n_6674 ^ mul_34_17_n_6677);
 assign mul_34_17_n_7188 = ~(mul_34_17_n_6673 ^ mul_34_17_n_94);
 assign mul_34_17_n_7187 = ~(mul_34_17_n_82 ^ mul_34_17_n_6594);
 assign mul_34_17_n_7186 = (mul_34_17_n_6667 ^ mul_34_17_n_6270);
 assign mul_34_17_n_7185 = ~(mul_34_17_n_11515 ^ mul_34_17_n_11516);
 assign mul_34_17_n_7388 = ~(mul_34_17_n_6402 ^ mul_34_17_n_6682);
 assign mul_34_17_n_7184 = (mul_34_17_n_11514 ^ mul_34_17_n_1);
 assign mul_34_17_n_7183 = ~(mul_34_17_n_5469 ^ (mul_34_17_n_4736 ^ (mul_34_17_n_5177 ^ mul_34_17_n_4726)));
 assign mul_34_17_n_7182 = (mul_34_17_n_83 ^ mul_34_17_n_84);
 assign mul_34_17_n_7181 = (mul_34_17_n_144 ^ mul_34_17_n_143);
 assign mul_34_17_n_7387 = ~(mul_34_17_n_5488 ^ (mul_34_17_n_4812 ^ (mul_34_17_n_5489 ^ mul_34_17_n_4116)));
 assign mul_34_17_n_7386 = ~(mul_34_17_n_5491 ^ (mul_34_17_n_3095 ^ (mul_34_17_n_5490 ^ mul_34_17_n_4468)));
 assign mul_34_17_n_7180 = ~(mul_34_17_n_6661 ^ mul_34_17_n_28);
 assign mul_34_17_n_7179 = ~(mul_34_17_n_139 ^ (mul_34_17_n_4065 ^ (mul_34_17_n_5471 ^ mul_34_17_n_3085)));
 assign mul_34_17_n_7178 = (mul_34_17_n_5551 ^ mul_34_17_n_6611);
 assign mul_34_17_n_7385 = ((mul_34_17_n_5540 & mul_34_17_n_5778) | ((mul_34_17_n_5540 & mul_34_17_n_5114)
    | (mul_34_17_n_5114 & mul_34_17_n_5778)));
 assign mul_34_17_n_7384 = ((mul_34_17_n_6115 & mul_34_17_n_4875) | ((mul_34_17_n_6115 & mul_34_17_n_2867)
    | (mul_34_17_n_2867 & mul_34_17_n_4875)));
 assign mul_34_17_n_7177 = (mul_34_17_n_6614 ^ mul_34_17_n_6610);
 assign mul_34_17_n_7176 = ~(mul_34_17_n_5457 ^ (mul_34_17_n_4181 ^ (mul_34_17_n_5458 ^ mul_34_17_n_2853)));
 assign mul_34_17_n_7175 = (mul_34_17_n_15 ^ mul_34_17_n_16);
 assign mul_34_17_n_7174 = ~(mul_34_17_n_5152 ^ (mul_34_17_n_3716 ^ (mul_34_17_n_4837 ^ mul_34_17_n_4680)));
 assign mul_34_17_n_7173 = (mul_34_17_n_115 ^ mul_34_17_n_6564);
 assign mul_34_17_n_7383 = ((mul_34_17_n_5693 & mul_34_17_n_5518) | ((mul_34_17_n_5693 & mul_34_17_n_5765)
    | (mul_34_17_n_5765 & mul_34_17_n_5518)));
 assign mul_34_17_n_7172 = (mul_34_17_n_6540 ^ mul_34_17_n_6535);
 assign mul_34_17_n_7171 = (mul_34_17_n_6590 ^ mul_34_17_n_6589);
 assign mul_34_17_n_7170 = (mul_34_17_n_58 ^ mul_34_17_n_6585);
 assign mul_34_17_n_7169 = ~(mul_34_17_n_5460 ^ (mul_34_17_n_4664 ^ (mul_34_17_n_5459 ^ mul_34_17_n_3824)));
 assign mul_34_17_n_7168 = (mul_34_17_n_6593 ^ mul_34_17_n_6648);
 assign mul_34_17_n_7167 = (mul_34_17_n_6663 ^ mul_34_17_n_6529);
 assign mul_34_17_n_7166 = (mul_34_17_n_6602 ^ mul_34_17_n_6601);
 assign mul_34_17_n_7382 = ((mul_34_17_n_5567 & mul_34_17_n_5725) | ((mul_34_17_n_5567 & mul_34_17_n_5675)
    | (mul_34_17_n_5675 & mul_34_17_n_5725)));
 assign mul_34_17_n_7381 = ((mul_34_17_n_6015 & mul_34_17_n_6678) | ((mul_34_17_n_6015 & mul_34_17_n_6016)
    | (mul_34_17_n_6016 & mul_34_17_n_6678)));
 assign mul_34_17_n_7380 = ((mul_34_17_n_5659 & mul_34_17_n_5796) | ((mul_34_17_n_5659 & mul_34_17_n_5715)
    | (mul_34_17_n_5715 & mul_34_17_n_5796)));
 assign mul_34_17_n_7379 = ((mul_34_17_n_5805 & mul_34_17_n_6680) | ((mul_34_17_n_5805 & mul_34_17_n_5804)
    | (mul_34_17_n_5804 & mul_34_17_n_6680)));
 assign mul_34_17_n_7378 = ((mul_34_17_n_5605 & mul_34_17_n_61) | ((mul_34_17_n_5605 & mul_34_17_n_5606)
    | (mul_34_17_n_5606 & mul_34_17_n_61)));
 assign mul_34_17_n_7377 = ((mul_34_17_n_5607 & mul_34_17_n_137) | ((mul_34_17_n_5607 & mul_34_17_n_6005)
    | (mul_34_17_n_6005 & mul_34_17_n_137)));
 assign mul_34_17_n_7376 = ((mul_34_17_n_5711 & mul_34_17_n_5773) | ((mul_34_17_n_5711 & mul_34_17_n_5712)
    | (mul_34_17_n_5712 & mul_34_17_n_5773)));
 assign mul_34_17_n_7375 = ((mul_34_17_n_5544 & mul_34_17_n_5720) | ((mul_34_17_n_5544 & mul_34_17_n_5542)
    | (mul_34_17_n_5542 & mul_34_17_n_5720)));
 assign mul_34_17_n_7374 = ((mul_34_17_n_5945 & mul_34_17_n_6010) | ((mul_34_17_n_5945 & mul_34_17_n_5887)
    | (mul_34_17_n_5887 & mul_34_17_n_6010)));
 assign mul_34_17_n_7373 = ((mul_34_17_n_5888 & mul_34_17_n_6368) | ((mul_34_17_n_5888 & mul_34_17_n_4896)
    | (mul_34_17_n_4896 & mul_34_17_n_6368)));
 assign mul_34_17_n_7372 = ((mul_34_17_n_5973 & mul_34_17_n_6048) | ((mul_34_17_n_5973 & mul_34_17_n_4412)
    | (mul_34_17_n_4412 & mul_34_17_n_6048)));
 assign mul_34_17_n_7371 = ((mul_34_17_n_5636 & mul_34_17_n_5791) | ((mul_34_17_n_5636 & mul_34_17_n_5637)
    | (mul_34_17_n_5637 & mul_34_17_n_5791)));
 assign mul_34_17_n_7370 = ((mul_34_17_n_5978 & mul_34_17_n_6107) | ((mul_34_17_n_5978 & mul_34_17_n_5976)
    | (mul_34_17_n_5976 & mul_34_17_n_6107)));
 assign mul_34_17_n_7368 = ((mul_34_17_n_5676 & mul_34_17_n_5762) | ((mul_34_17_n_5676 & mul_34_17_n_5680)
    | (mul_34_17_n_5680 & mul_34_17_n_5762)));
 assign mul_34_17_n_7367 = ((mul_34_17_n_5679 & mul_34_17_n_6080) | ((mul_34_17_n_5679 & mul_34_17_n_6007)
    | (mul_34_17_n_6007 & mul_34_17_n_6080)));
 assign mul_34_17_n_7365 = ((mul_34_17_n_4903 & mul_34_17_n_3004) | (mul_34_17_n_6442 & mul_34_17_n_6436));
 assign mul_34_17_n_7364 = ((mul_34_17_n_5709 & mul_34_17_n_5770) | ((mul_34_17_n_5709 & mul_34_17_n_5120)
    | (mul_34_17_n_5120 & mul_34_17_n_5770)));
 assign mul_34_17_n_7363 = ((mul_34_17_n_5561 & mul_34_17_n_5799) | ((mul_34_17_n_5561 & mul_34_17_n_5537)
    | (mul_34_17_n_5537 & mul_34_17_n_5799)));
 assign mul_34_17_n_7362 = ((mul_34_17_n_113 & mul_34_17_n_5741) | ((mul_34_17_n_113 & mul_34_17_n_49)
    | (mul_34_17_n_49 & mul_34_17_n_5741)));
 assign mul_34_17_n_7361 = ((mul_34_17_n_5543 & mul_34_17_n_5777) | ((mul_34_17_n_5543 & mul_34_17_n_5545)
    | (mul_34_17_n_5545 & mul_34_17_n_5777)));
 assign mul_34_17_n_7360 = ((mul_34_17_n_5514 & mul_34_17_n_5775) | ((mul_34_17_n_5514 & mul_34_17_n_5536)
    | (mul_34_17_n_5536 & mul_34_17_n_5775)));
 assign mul_34_17_n_7359 = ((mul_34_17_n_5970 & mul_34_17_n_6062) | ((mul_34_17_n_5970 & mul_34_17_n_5969)
    | (mul_34_17_n_5969 & mul_34_17_n_6062)));
 assign mul_34_17_n_7358 = ((mul_34_17_n_5997 & mul_34_17_n_6075) | ((mul_34_17_n_5997 & mul_34_17_n_5995)
    | (mul_34_17_n_5995 & mul_34_17_n_6075)));
 assign mul_34_17_n_7356 = ((mul_34_17_n_6032 & mul_34_17_n_6093) | ((mul_34_17_n_6032 & mul_34_17_n_5941)
    | (mul_34_17_n_5941 & mul_34_17_n_6093)));
 assign mul_34_17_n_7355 = ((mul_34_17_n_6014 & mul_34_17_n_6085) | ((mul_34_17_n_6014 & mul_34_17_n_5638)
    | (mul_34_17_n_5638 & mul_34_17_n_6085)));
 assign mul_34_17_n_7354 = ((mul_34_17_n_5701 & mul_34_17_n_5768) | ((mul_34_17_n_5701 & mul_34_17_n_5700)
    | (mul_34_17_n_5700 & mul_34_17_n_5768)));
 assign mul_34_17_n_7353 = ((mul_34_17_n_131 & mul_34_17_n_129) | ((mul_34_17_n_131 & mul_34_17_n_133)
    | (mul_34_17_n_133 & mul_34_17_n_129)));
 assign mul_34_17_n_7352 = ((mul_34_17_n_5965 & mul_34_17_n_5695) | ((mul_34_17_n_5965 & mul_34_17_n_5981)
    | (mul_34_17_n_5981 & mul_34_17_n_5695)));
 assign mul_34_17_n_7351 = ((mul_34_17_n_5425 & mul_34_17_n_6665) | ((mul_34_17_n_5425 & mul_34_17_n_108)
    | (mul_34_17_n_108 & mul_34_17_n_6665)));
 assign mul_34_17_n_7350 = ((mul_34_17_n_6036 & mul_34_17_n_6633) | ((mul_34_17_n_6036 & mul_34_17_n_5891)
    | (mul_34_17_n_5891 & mul_34_17_n_6633)));
 assign mul_34_17_n_7347 = ((mul_34_17_n_6028 & mul_34_17_n_6094) | ((mul_34_17_n_6028 & mul_34_17_n_6026)
    | (mul_34_17_n_6026 & mul_34_17_n_6094)));
 assign mul_34_17_n_7346 = ((mul_34_17_n_5667 & mul_34_17_n_6400) | ((mul_34_17_n_5667 & mul_34_17_n_5671)
    | (mul_34_17_n_5671 & mul_34_17_n_6400)));
 assign mul_34_17_n_7345 = ((mul_34_17_n_5697 & mul_34_17_n_5766) | ((mul_34_17_n_5697 & mul_34_17_n_5691)
    | (mul_34_17_n_5691 & mul_34_17_n_5766)));
 assign mul_34_17_n_7344 = ((mul_34_17_n_5999 & mul_34_17_n_6105) | ((mul_34_17_n_5999 & mul_34_17_n_6013)
    | (mul_34_17_n_6013 & mul_34_17_n_6105)));
 assign mul_34_17_n_7343 = ((mul_34_17_n_5656 & mul_34_17_n_6079) | ((mul_34_17_n_5656 & mul_34_17_n_3033)
    | (mul_34_17_n_3033 & mul_34_17_n_6079)));
 assign mul_34_17_n_7342 = ((mul_34_17_n_5534 & mul_34_17_n_5752) | ((mul_34_17_n_5534 & mul_34_17_n_4887)
    | (mul_34_17_n_4887 & mul_34_17_n_5752)));
 assign mul_34_17_n_7341 = ((mul_34_17_n_6027 & mul_34_17_n_6040) | ((mul_34_17_n_6027 & mul_34_17_n_6030)
    | (mul_34_17_n_6030 & mul_34_17_n_6040)));
 assign mul_34_17_n_7340 = ((mul_34_17_n_5966 & mul_34_17_n_6061) | ((mul_34_17_n_5966 & mul_34_17_n_3023)
    | (mul_34_17_n_3023 & mul_34_17_n_6061)));
 assign mul_34_17_n_7339 = ((mul_34_17_n_5525 & mul_34_17_n_6361) | ((mul_34_17_n_5525 & mul_34_17_n_5661)
    | (mul_34_17_n_5661 & mul_34_17_n_6361)));
 assign mul_34_17_n_7338 = ((mul_34_17_n_5584 & mul_34_17_n_6042) | ((mul_34_17_n_5584 & mul_34_17_n_4895)
    | (mul_34_17_n_4895 & mul_34_17_n_6042)));
 assign mul_34_17_n_7337 = ((mul_34_17_n_5685 & mul_34_17_n_6087) | ((mul_34_17_n_5685 & mul_34_17_n_4892)
    | (mul_34_17_n_4892 & mul_34_17_n_6087)));
 assign mul_34_17_n_7336 = ((mul_34_17_n_5554 & mul_34_17_n_6389) | ((mul_34_17_n_5554 & mul_34_17_n_5112)
    | (mul_34_17_n_5112 & mul_34_17_n_6389)));
 assign mul_34_17_n_7335 = ((mul_34_17_n_5684 & mul_34_17_n_6086) | ((mul_34_17_n_5684 & mul_34_17_n_6017)
    | (mul_34_17_n_6017 & mul_34_17_n_6086)));
 assign mul_34_17_n_7334 = ((mul_34_17_n_6002 & mul_34_17_n_6077) | ((mul_34_17_n_6002 & mul_34_17_n_4898)
    | (mul_34_17_n_4898 & mul_34_17_n_6077)));
 assign mul_34_17_n_7333 = ((mul_34_17_n_5682 & mul_34_17_n_6083) | ((mul_34_17_n_5682 & mul_34_17_n_5899)
    | (mul_34_17_n_5899 & mul_34_17_n_6083)));
 assign mul_34_17_n_7332 = ((mul_34_17_n_5683 & mul_34_17_n_6084) | ((mul_34_17_n_5683 & mul_34_17_n_6009)
    | (mul_34_17_n_6009 & mul_34_17_n_6084)));
 assign mul_34_17_n_7331 = ((mul_34_17_n_5907 & mul_34_17_n_6045) | ((mul_34_17_n_5907 & mul_34_17_n_5967)
    | (mul_34_17_n_5967 & mul_34_17_n_6045)));
 assign mul_34_17_n_7330 = ((mul_34_17_n_5205 & mul_34_17_n_6423) | ((mul_34_17_n_5205 & mul_34_17_n_5704)
    | (mul_34_17_n_5704 & mul_34_17_n_6423)));
 assign mul_34_17_n_7328 = ((mul_34_17_n_6020 & mul_34_17_n_6038) | ((mul_34_17_n_6020 & mul_34_17_n_3024)
    | (mul_34_17_n_3024 & mul_34_17_n_6038)));
 assign mul_34_17_n_7327 = ((mul_34_17_n_5977 & mul_34_17_n_6104) | ((mul_34_17_n_5977 & mul_34_17_n_4894)
    | (mul_34_17_n_4894 & mul_34_17_n_6104)));
 assign mul_34_17_n_7325 = ((mul_34_17_n_5624 & mul_34_17_n_5788) | ((mul_34_17_n_5624 & mul_34_17_n_5619)
    | (mul_34_17_n_5619 & mul_34_17_n_5788)));
 assign mul_34_17_n_7324 = ((mul_34_17_n_6035 & mul_34_17_n_6097) | ((mul_34_17_n_6035 & mul_34_17_n_5919)
    | (mul_34_17_n_5919 & mul_34_17_n_6097)));
 assign mul_34_17_n_7323 = ((mul_34_17_n_6037 & mul_34_17_n_6052) | ((mul_34_17_n_6037 & mul_34_17_n_4391)
    | (mul_34_17_n_4391 & mul_34_17_n_6052)));
 assign mul_34_17_n_7322 = ((mul_34_17_n_5666 & mul_34_17_n_5756) | ((mul_34_17_n_5666 & mul_34_17_n_5117)
    | (mul_34_17_n_5117 & mul_34_17_n_5756)));
 assign mul_34_17_n_7321 = ~(mul_34_17_n_11517 ^ mul_34_17_n_11518);
 assign mul_34_17_n_7320 = ((mul_34_17_n_5687 & mul_34_17_n_5740) | ((mul_34_17_n_5687 & mul_34_17_n_5692)
    | (mul_34_17_n_5692 & mul_34_17_n_5740)));
 assign mul_34_17_n_7318 = ((mul_34_17_n_5608 & mul_34_17_n_5737) | ((mul_34_17_n_5608 & mul_34_17_n_5109)
    | (mul_34_17_n_5109 & mul_34_17_n_5737)));
 assign mul_34_17_n_7317 = ((mul_34_17_n_5504 & mul_34_17_n_6098) | ((mul_34_17_n_5504 & mul_34_17_n_103)
    | (mul_34_17_n_103 & mul_34_17_n_6098)));
 assign mul_34_17_n_7315 = ((mul_34_17_n_5699 & mul_34_17_n_54) | ((mul_34_17_n_5699 & mul_34_17_n_5593)
    | (mul_34_17_n_5593 & mul_34_17_n_54)));
 assign mul_34_17_n_7314 = (mul_34_17_n_6607 ^ mul_34_17_n_6543);
 assign mul_34_17_n_7313 = ((mul_34_17_n_5927 & mul_34_17_n_6401) | ((mul_34_17_n_5927 & mul_34_17_n_5937)
    | (mul_34_17_n_5937 & mul_34_17_n_6401)));
 assign mul_34_17_n_7312 = ((mul_34_17_n_5558 & mul_34_17_n_147) | ((mul_34_17_n_5558 & mul_34_17_n_5942)
    | (mul_34_17_n_5942 & mul_34_17_n_147)));
 assign mul_34_17_n_7311 = ((mul_34_17_n_5943 & mul_34_17_n_6377) | ((mul_34_17_n_5943 & mul_34_17_n_5694)
    | (mul_34_17_n_5694 & mul_34_17_n_6377)));
 assign mul_34_17_n_7310 = ((mul_34_17_n_5642 & mul_34_17_n_5817) | (mul_34_17_n_6446 & mul_34_17_n_99));
 assign mul_34_17_n_7309 = ~((mul_34_17_n_5950 & mul_34_17_n_5953) | (mul_34_17_n_6388 & mul_34_17_n_6428));
 assign mul_34_17_n_7308 = ((mul_34_17_n_5917 & mul_34_17_n_6099) | ((mul_34_17_n_5917 & mul_34_17_n_5929)
    | (mul_34_17_n_5929 & mul_34_17_n_6099)));
 assign mul_34_17_n_7307 = ((mul_34_17_n_5616 & mul_34_17_n_5786) | ((mul_34_17_n_5616 & mul_34_17_n_5617)
    | (mul_34_17_n_5617 & mul_34_17_n_5786)));
 assign mul_34_17_n_7306 = (mul_34_17_n_31 ^ mul_34_17_n_29);
 assign mul_34_17_n_7305 = ((mul_34_17_n_6000 & mul_34_17_n_6106) | ((mul_34_17_n_6000 & mul_34_17_n_6006)
    | (mul_34_17_n_6006 & mul_34_17_n_6106)));
 assign mul_34_17_n_7304 = ((mul_34_17_n_5634 & mul_34_17_n_5748) | ((mul_34_17_n_5634 & mul_34_17_n_5690)
    | (mul_34_17_n_5690 & mul_34_17_n_5748)));
 assign mul_34_17_n_7303 = ~(mul_34_17_n_5486 ^ (mul_34_17_n_4717 ^ (mul_34_17_n_5485 ^ mul_34_17_n_4747)));
 assign mul_34_17_n_7302 = ((mul_34_17_n_5931 & mul_34_17_n_6688) | ((mul_34_17_n_5931 & mul_34_17_n_5933)
    | (mul_34_17_n_5933 & mul_34_17_n_6688)));
 assign mul_34_17_n_7301 = ((mul_34_17_n_5555 & mul_34_17_n_5774) | ((mul_34_17_n_5555 & mul_34_17_n_5580)
    | (mul_34_17_n_5580 & mul_34_17_n_5774)));
 assign mul_34_17_n_7299 = ((mul_34_17_n_5660 & mul_34_17_n_5757) | ((mul_34_17_n_5660 & mul_34_17_n_5601)
    | (mul_34_17_n_5601 & mul_34_17_n_5757)));
 assign mul_34_17_n_7298 = ((mul_34_17_n_5648 & mul_34_17_n_5742) | ((mul_34_17_n_5648 & mul_34_17_n_3962)
    | (mul_34_17_n_3962 & mul_34_17_n_5742)));
 assign mul_34_17_n_7297 = ((mul_34_17_n_5672 & mul_34_17_n_5761) | ((mul_34_17_n_5672 & mul_34_17_n_5670)
    | (mul_34_17_n_5670 & mul_34_17_n_5761)));
 assign mul_34_17_n_7296 = ~(mul_34_17_n_5470 ^ (mul_34_17_n_4687 ^ (mul_34_17_n_5472 ^ mul_34_17_n_4748)));
 assign mul_34_17_n_7295 = ((mul_34_17_n_5526 & mul_34_17_n_5801) | ((mul_34_17_n_5526 & mul_34_17_n_5535)
    | (mul_34_17_n_5535 & mul_34_17_n_5801)));
 assign mul_34_17_n_7293 = ((mul_34_17_n_5589 & mul_34_17_n_6103) | ((mul_34_17_n_5589 & mul_34_17_n_5955)
    | (mul_34_17_n_5955 & mul_34_17_n_6103)));
 assign mul_34_17_n_7292 = ((mul_34_17_n_5513 & mul_34_17_n_5780) | ((mul_34_17_n_5513 & mul_34_17_n_3961)
    | (mul_34_17_n_3961 & mul_34_17_n_5780)));
 assign mul_34_17_n_7291 = ((mul_34_17_n_5538 & mul_34_17_n_5717) | ((mul_34_17_n_5538 & mul_34_17_n_5662)
    | (mul_34_17_n_5662 & mul_34_17_n_5717)));
 assign mul_34_17_n_7290 = ((mul_34_17_n_6031 & mul_34_17_n_6095) | ((mul_34_17_n_6031 & mul_34_17_n_5429)
    | (mul_34_17_n_5429 & mul_34_17_n_6095)));
 assign mul_34_17_n_7165 = ~mul_34_17_n_7044;
 assign mul_34_17_n_7163 = ~mul_34_17_n_7162;
 assign mul_34_17_n_7161 = ~mul_34_17_n_7160;
 assign mul_34_17_n_7151 = ~mul_34_17_n_7150;
 assign mul_34_17_n_7134 = ~mul_34_17_n_7133;
 assign mul_34_17_n_7131 = ~mul_34_17_n_7130;
 assign mul_34_17_n_7127 = ~mul_34_17_n_7126;
 assign mul_34_17_n_7122 = ~mul_34_17_n_7121;
 assign mul_34_17_n_7107 = ~mul_34_17_n_7106;
 assign mul_34_17_n_7102 = ~mul_34_17_n_7103;
 assign mul_34_17_n_7096 = ~mul_34_17_n_7095;
 assign mul_34_17_n_7083 = ~mul_34_17_n_7082;
 assign mul_34_17_n_7063 = ~mul_34_17_n_7062;
 assign mul_34_17_n_7060 = ~mul_34_17_n_7059;
 assign mul_34_17_n_7054 = ~mul_34_17_n_7055;
 assign mul_34_17_n_7053 = ~mul_34_17_n_7052;
 assign mul_34_17_n_7048 = ~(mul_34_17_n_5143 ^ (mul_34_17_n_4857 ^ (mul_34_17_n_5189 ^ mul_34_17_n_3670)));
 assign mul_34_17_n_7046 = ~(mul_34_17_n_5463 ^ (mul_34_17_n_3391 ^ (mul_34_17_n_5478 ^ mul_34_17_n_3115)));
 assign mul_34_17_n_7044 = ((mul_34_17_n_5693 & mul_34_17_n_5765) | ((mul_34_17_n_5693 & mul_34_17_n_5518)
    | (mul_34_17_n_5518 & mul_34_17_n_5765)));
 assign mul_34_17_n_7043 = (mul_34_17_n_6218 ^ mul_34_17_n_6182);
 assign mul_34_17_n_7038 = ~(mul_34_17_n_5146 ^ (mul_34_17_n_3697 ^ (mul_34_17_n_5147 ^ mul_34_17_n_3138)));
 assign mul_34_17_n_7028 = ~(mul_34_17_n_5161 ^ (mul_34_17_n_3787 ^ (mul_34_17_n_5159 ^ mul_34_17_n_3767)));
 assign mul_34_17_n_7027 = (mul_34_17_n_6166 ^ mul_34_17_n_6209);
 assign mul_34_17_n_7024 = ~(mul_34_17_n_5182 ^ (mul_34_17_n_3900 ^ (mul_34_17_n_5183 ^ mul_34_17_n_4695)));
 assign mul_34_17_n_7022 = ~(mul_34_17_n_6171 ^ mul_34_17_n_6212);
 assign mul_34_17_n_7020 = ~(mul_34_17_n_6183 ^ mul_34_17_n_6177);
 assign mul_34_17_n_7019 = ~(mul_34_17_n_5195 ^ (mul_34_17_n_3850 ^ (mul_34_17_n_5196 ^ mul_34_17_n_3722)));
 assign mul_34_17_n_7014 = (mul_34_17_n_6168 ^ mul_34_17_n_6202);
 assign mul_34_17_n_7012 = ~(mul_34_17_n_6198 ^ mul_34_17_n_5411);
 assign mul_34_17_n_7011 = ~(mul_34_17_n_5168 ^ (mul_34_17_n_3805 ^ (mul_34_17_n_5194 ^ mul_34_17_n_3920)));
 assign mul_34_17_n_7002 = ~(mul_34_17_n_6504 ^ mul_34_17_n_136);
 assign mul_34_17_n_7000 = ~(mul_34_17_n_5160 ^ (mul_34_17_n_3770 ^ (mul_34_17_n_5162 ^ mul_34_17_n_3418)));
 assign mul_34_17_n_6995 = (mul_34_17_n_6208 ^ mul_34_17_n_6165);
 assign mul_34_17_n_6994 = ~(mul_34_17_n_6197 ^ mul_34_17_n_6169);
 assign mul_34_17_n_6993 = ~(mul_34_17_n_5179 ^ (mul_34_17_n_3846 ^ (mul_34_17_n_5181 ^ mul_34_17_n_4690)));
 assign mul_34_17_n_6992 = ~(mul_34_17_n_5482 ^ (mul_34_17_n_3745 ^ (mul_34_17_n_5178 ^ mul_34_17_n_3686)));
 assign mul_34_17_n_6990 = ~(mul_34_17_n_6179 ^ mul_34_17_n_6213);
 assign mul_34_17_n_6989 = ~(mul_34_17_n_5190 ^ (mul_34_17_n_3552 ^ (mul_34_17_n_5188 ^ mul_34_17_n_3731)));
 assign mul_34_17_n_6987 = ~(mul_34_17_n_6155 ^ mul_34_17_n_4907);
 assign mul_34_17_n_6985 = ~(mul_34_17_n_5200 ^ (mul_34_17_n_4604 ^ (mul_34_17_n_5184 ^ mul_34_17_n_3886)));
 assign mul_34_17_n_6984 = ((mul_34_17_n_3660 | mul_34_17_n_3064) & (mul_34_17_n_6155 | mul_34_17_n_6356));
 assign mul_34_17_n_6983 = ~(mul_34_17_n_5164 ^ (mul_34_17_n_3780 ^ (mul_34_17_n_5163 ^ mul_34_17_n_3777)));
 assign mul_34_17_n_6979 = ~(mul_34_17_n_5174 ^ (mul_34_17_n_3897 ^ (mul_34_17_n_5496 ^ mul_34_17_n_3615)));
 assign mul_34_17_n_6978 = (mul_34_17_n_6167 ^ mul_34_17_n_6196);
 assign mul_34_17_n_6976 = ~(mul_34_17_n_6334 ^ mul_34_17_n_6546);
 assign mul_34_17_n_6975 = ~(mul_34_17_n_6517 ^ mul_34_17_n_6487);
 assign mul_34_17_n_6974 = ~(mul_34_17_n_5493 ^ (mul_34_17_n_4187 ^ (mul_34_17_n_5468 ^ mul_34_17_n_4246)));
 assign mul_34_17_n_6971 = ((mul_34_17_n_5137 | mul_34_17_n_3062) & (mul_34_17_n_6188 | mul_34_17_n_6295));
 assign mul_34_17_n_6970 = ~(mul_34_17_n_5158 ^ (mul_34_17_n_3296 ^ (mul_34_17_n_5197 ^ mul_34_17_n_3828)));
 assign mul_34_17_n_6969 = ~(mul_34_17_n_5154 ^ (mul_34_17_n_4659 ^ (mul_34_17_n_3660 ^ mul_34_17_n_3064)));
 assign mul_34_17_n_6967 = ~(mul_34_17_n_6159 ^ mul_34_17_n_6211);
 assign mul_34_17_n_7164 = ((mul_34_17_n_6308 & mul_34_17_n_5108) | (mul_34_17_n_6307 & mul_34_17_n_5987));
 assign mul_34_17_n_6966 = (mul_34_17_n_64 ^ mul_34_17_n_6609);
 assign mul_34_17_n_6965 = (mul_34_17_n_35 ^ mul_34_17_n_36);
 assign mul_34_17_n_6964 = (mul_34_17_n_6399 ^ mul_34_17_n_6228);
 assign mul_34_17_n_7162 = (mul_34_17_n_5987 ^ mul_34_17_n_6307);
 assign mul_34_17_n_7160 = ~(mul_34_17_n_6309 ^ mul_34_17_n_5108);
 assign mul_34_17_n_6963 = ~(mul_34_17_n_5473 ^ (mul_34_17_n_4602 ^ (mul_34_17_n_5498 ^ mul_34_17_n_3028)));
 assign mul_34_17_n_7159 = ~(mul_34_17_n_6305 ^ mul_34_17_n_6676);
 assign mul_34_17_n_6962 = (mul_34_17_n_5595 ^ mul_34_17_n_6318);
 assign mul_34_17_n_6961 = ~(mul_34_17_n_5165 ^ (mul_34_17_n_3823 ^ (mul_34_17_n_3934 ^ mul_34_17_n_3746)));
 assign mul_34_17_n_6960 = (mul_34_17_n_6379 ^ mul_34_17_n_6283);
 assign mul_34_17_n_6959 = (mul_34_17_n_6357 ^ mul_34_17_n_6324);
 assign mul_34_17_n_6958 = (mul_34_17_n_6224 ^ mul_34_17_n_6226);
 assign mul_34_17_n_6957 = ~(mul_34_17_n_5201 ^ (mul_34_17_n_3848 ^ (mul_34_17_n_3937 ^ mul_34_17_n_3815)));
 assign mul_34_17_n_6956 = ~(mul_34_17_n_4870 ^ (mul_34_17_n_5454 ^ (mul_34_17_n_5187 ^ mul_34_17_n_3879)));
 assign mul_34_17_n_6955 = (mul_34_17_n_6260 ^ mul_34_17_n_21);
 assign mul_34_17_n_6954 = (mul_34_17_n_37 ^ mul_34_17_n_6277);
 assign mul_34_17_n_6953 = (mul_34_17_n_6242 ^ mul_34_17_n_6241);
 assign mul_34_17_n_6952 = (mul_34_17_n_6239 ^ mul_34_17_n_6323);
 assign mul_34_17_n_6951 = ~(mul_34_17_n_5171 ^ (mul_34_17_n_4865 ^ (mul_34_17_n_5199 ^ mul_34_17_n_3587)));
 assign mul_34_17_n_6950 = ~(mul_34_17_n_6364 ^ mul_34_17_n_5136);
 assign mul_34_17_n_6949 = (mul_34_17_n_6236 ^ mul_34_17_n_5714);
 assign mul_34_17_n_6948 = (mul_34_17_n_6375 ^ mul_34_17_n_6227);
 assign mul_34_17_n_6947 = (mul_34_17_n_5118 ^ mul_34_17_n_6249);
 assign mul_34_17_n_7158 = ~(mul_34_17_n_4864 ^ (mul_34_17_n_5149 ^ (mul_34_17_n_5151 ^ mul_34_17_n_3715)));
 assign mul_34_17_n_6946 = (mul_34_17_n_6225 ^ mul_34_17_n_10);
 assign mul_34_17_n_6945 = ~(mul_34_17_n_5150 ^ (mul_34_17_n_3208 ^ (mul_34_17_n_5148 ^ mul_34_17_n_4571)));
 assign mul_34_17_n_6944 = (mul_34_17_n_6618 ^ mul_34_17_n_6552);
 assign mul_34_17_n_6943 = (mul_34_17_n_6278 ^ mul_34_17_n_6630);
 assign mul_34_17_n_7157 = (mul_34_17_n_6235 ^ mul_34_17_n_5140);
 assign mul_34_17_n_6942 = (mul_34_17_n_93 ^ mul_34_17_n_6574);
 assign mul_34_17_n_6941 = ~(mul_34_17_n_5475 ^ (mul_34_17_n_4589 ^ (mul_34_17_n_5476 ^ mul_34_17_n_3532)));
 assign mul_34_17_n_6940 = (mul_34_17_n_6394 ^ mul_34_17_n_6246);
 assign mul_34_17_n_6939 = (mul_34_17_n_6255 ^ mul_34_17_n_6250);
 assign mul_34_17_n_6938 = (mul_34_17_n_6586 ^ mul_34_17_n_6627);
 assign mul_34_17_n_6937 = ~(mul_34_17_n_91 ^ mul_34_17_n_81);
 assign mul_34_17_n_7156 = ((mul_34_17_n_5135 & mul_34_17_n_6364) | ((mul_34_17_n_5135 & mul_34_17_n_5898)
    | (mul_34_17_n_5898 & mul_34_17_n_6364)));
 assign mul_34_17_n_7155 = ((mul_34_17_n_5119 & mul_34_17_n_5885) | ((mul_34_17_n_5119 & mul_34_17_n_5505)
    | (mul_34_17_n_5505 & mul_34_17_n_5885)));
 assign mul_34_17_n_7154 = ((mul_34_17_n_5713 & mul_34_17_n_6043) | ((mul_34_17_n_5713 & mul_34_17_n_6024)
    | (mul_34_17_n_6024 & mul_34_17_n_6043)));
 assign mul_34_17_n_7153 = ((mul_34_17_n_5629 & mul_34_17_n_6217) | ((mul_34_17_n_5629 & mul_34_17_n_5627)
    | (mul_34_17_n_5627 & mul_34_17_n_6217)));
 assign mul_34_17_n_7152 = ((mul_34_17_n_5644 & mul_34_17_n_5745) | ((mul_34_17_n_5644 & mul_34_17_n_5626)
    | (mul_34_17_n_5626 & mul_34_17_n_5745)));
 assign mul_34_17_n_7150 = ((mul_34_17_n_5956 & mul_34_17_n_5782) | ((mul_34_17_n_5956 & mul_34_17_n_5959)
    | (mul_34_17_n_5959 & mul_34_17_n_5782)));
 assign mul_34_17_n_7149 = ((mul_34_17_n_6022 & mul_34_17_n_6090) | ((mul_34_17_n_6022 & mul_34_17_n_6023)
    | (mul_34_17_n_6023 & mul_34_17_n_6090)));
 assign mul_34_17_n_7148 = ~(mul_34_17_n_6146 ^ mul_34_17_n_5688);
 assign mul_34_17_n_7147 = ((mul_34_17_n_5643 & mul_34_17_n_5750) | ((mul_34_17_n_5643 & mul_34_17_n_5579)
    | (mul_34_17_n_5579 & mul_34_17_n_5750)));
 assign mul_34_17_n_7146 = ~(mul_34_17_n_6429 ^ mul_34_17_n_5872);
 assign mul_34_17_n_7145 = ((mul_34_17_n_5890 & mul_34_17_n_85) | ((mul_34_17_n_5890 & mul_34_17_n_5615)
    | (mul_34_17_n_5615 & mul_34_17_n_85)));
 assign mul_34_17_n_7144 = ((mul_34_17_n_5610 & mul_34_17_n_5738) | ((mul_34_17_n_5610 & mul_34_17_n_5926)
    | (mul_34_17_n_5926 & mul_34_17_n_5738)));
 assign mul_34_17_n_7143 = ((mul_34_17_n_5633 & mul_34_17_n_105) | ((mul_34_17_n_5633 & mul_34_17_n_5628)
    | (mul_34_17_n_5628 & mul_34_17_n_105)));
 assign mul_34_17_n_7142 = ((mul_34_17_n_5651 & mul_34_17_n_5753) | ((mul_34_17_n_5651 & mul_34_17_n_6033)
    | (mul_34_17_n_6033 & mul_34_17_n_5753)));
 assign mul_34_17_n_7141 = ((mul_34_17_n_5522 & mul_34_17_n_5716) | ((mul_34_17_n_5522 & mul_34_17_n_5653)
    | (mul_34_17_n_5653 & mul_34_17_n_5716)));
 assign mul_34_17_n_7140 = ((mul_34_17_n_5895 & mul_34_17_n_5792) | ((mul_34_17_n_5895 & mul_34_17_n_5904)
    | (mul_34_17_n_5904 & mul_34_17_n_5792)));
 assign mul_34_17_n_7139 = ((mul_34_17_n_5975 & mul_34_17_n_5783) | ((mul_34_17_n_5975 & mul_34_17_n_5971)
    | (mul_34_17_n_5971 & mul_34_17_n_5783)));
 assign mul_34_17_n_7138 = ((mul_34_17_n_5647 & mul_34_17_n_5751) | ((mul_34_17_n_5647 & mul_34_17_n_5646)
    | (mul_34_17_n_5646 & mul_34_17_n_5751)));
 assign mul_34_17_n_7137 = ((mul_34_17_n_5602 & mul_34_17_n_5754) | ((mul_34_17_n_5602 & mul_34_17_n_5639)
    | (mul_34_17_n_5639 & mul_34_17_n_5754)));
 assign mul_34_17_n_7136 = ((mul_34_17_n_5900 & mul_34_17_n_6049) | ((mul_34_17_n_5900 & mul_34_17_n_5908)
    | (mul_34_17_n_5908 & mul_34_17_n_6049)));
 assign mul_34_17_n_7135 = ~(mul_34_17_n_6147 ^ mul_34_17_n_5577);
 assign mul_34_17_n_7133 = ((mul_34_17_n_5564 & mul_34_17_n_5724) | ((mul_34_17_n_5564 & mul_34_17_n_5566)
    | (mul_34_17_n_5566 & mul_34_17_n_5724)));
 assign mul_34_17_n_7132 = ((mul_34_17_n_5960 & mul_34_17_n_6041) | ((mul_34_17_n_5960 & mul_34_17_n_5910)
    | (mul_34_17_n_5910 & mul_34_17_n_6041)));
 assign mul_34_17_n_7130 = ((mul_34_17_n_5552 & mul_34_17_n_5722) | ((mul_34_17_n_5552 & mul_34_17_n_5553)
    | (mul_34_17_n_5553 & mul_34_17_n_5722)));
 assign mul_34_17_n_7129 = ((mul_34_17_n_56 & mul_34_17_n_5803) | ((mul_34_17_n_56 & mul_34_17_n_5609)
    | (mul_34_17_n_5609 & mul_34_17_n_5803)));
 assign mul_34_17_n_7128 = ((mul_34_17_n_5592 & mul_34_17_n_5731) | ((mul_34_17_n_5592 & mul_34_17_n_5594)
    | (mul_34_17_n_5594 & mul_34_17_n_5731)));
 assign mul_34_17_n_7126 = ((mul_34_17_n_5658 & mul_34_17_n_5793) | ((mul_34_17_n_5658 & mul_34_17_n_5621)
    | (mul_34_17_n_5621 & mul_34_17_n_5793)));
 assign mul_34_17_n_7125 = ((mul_34_17_n_5570 & mul_34_17_n_5795) | ((mul_34_17_n_5570 & mul_34_17_n_5571)
    | (mul_34_17_n_5571 & mul_34_17_n_5795)));
 assign mul_34_17_n_7124 = ((mul_34_17_n_5688 & mul_34_17_n_5447) | ((mul_34_17_n_5688 & mul_34_17_n_4040)
    | (mul_34_17_n_4040 & mul_34_17_n_5447)));
 assign mul_34_17_n_7123 = ((mul_34_17_n_5650 & mul_34_17_n_5449) | ((mul_34_17_n_5650 & mul_34_17_n_5652)
    | (mul_34_17_n_5652 & mul_34_17_n_5449)));
 assign mul_34_17_n_7121 = ((mul_34_17_n_75 & mul_34_17_n_6053) | ((mul_34_17_n_75 & mul_34_17_n_5946)
    | (mul_34_17_n_5946 & mul_34_17_n_6053)));
 assign mul_34_17_n_7120 = ((mul_34_17_n_5948 & mul_34_17_n_6057) | ((mul_34_17_n_5948 & mul_34_17_n_5905)
    | (mul_34_17_n_5905 & mul_34_17_n_6057)));
 assign mul_34_17_n_7119 = ((mul_34_17_n_4905 & mul_34_17_n_6138) | ((mul_34_17_n_4905 & mul_34_17_n_5923)
    | (mul_34_17_n_5923 & mul_34_17_n_6138)));
 assign mul_34_17_n_7118 = ((mul_34_17_n_5954 & mul_34_17_n_6055) | ((mul_34_17_n_5954 & mul_34_17_n_5957)
    | (mul_34_17_n_5957 & mul_34_17_n_6055)));
 assign mul_34_17_n_7117 = (mul_34_17_n_6360 ^ mul_34_17_n_6336);
 assign mul_34_17_n_6936 = ~(mul_34_17_n_5497 ^ (mul_34_17_n_4574 ^ (mul_34_17_n_5176 ^ mul_34_17_n_4572)));
 assign mul_34_17_n_7116 = ((mul_34_17_n_5962 & mul_34_17_n_6058) | ((mul_34_17_n_5962 & mul_34_17_n_5963)
    | (mul_34_17_n_5963 & mul_34_17_n_6058)));
 assign mul_34_17_n_7115 = ((mul_34_17_n_5875 & mul_34_17_n_6056) | ((mul_34_17_n_5875 & mul_34_17_n_5916)
    | (mul_34_17_n_5916 & mul_34_17_n_6056)));
 assign mul_34_17_n_7114 = ((mul_34_17_n_5596 & mul_34_17_n_5760) | ((mul_34_17_n_5596 & mul_34_17_n_5541)
    | (mul_34_17_n_5541 & mul_34_17_n_5760)));
 assign mul_34_17_n_7113 = ((mul_34_17_n_5631 & mul_34_17_n_5771) | ((mul_34_17_n_5631 & mul_34_17_n_5588)
    | (mul_34_17_n_5588 & mul_34_17_n_5771)));
 assign mul_34_17_n_7112 = (mul_34_17_n_39 ^ mul_34_17_n_40);
 assign mul_34_17_n_7111 = (mul_34_17_n_6369 ^ mul_34_17_n_6286);
 assign mul_34_17_n_7110 = (mul_34_17_n_6335 ^ mul_34_17_n_6333);
 assign mul_34_17_n_7109 = ((mul_34_17_n_5107 & mul_34_17_n_5744) | ((mul_34_17_n_5107 & mul_34_17_n_5625)
    | (mul_34_17_n_5625 & mul_34_17_n_5744)));
 assign mul_34_17_n_7108 = ~(mul_34_17_n_5166 ^ (mul_34_17_n_4001 ^ (mul_34_17_n_5167 ^ mul_34_17_n_4339)));
 assign mul_34_17_n_7106 = ((mul_34_17_n_5597 & mul_34_17_n_6069) | ((mul_34_17_n_5597 & mul_34_17_n_5980)
    | (mul_34_17_n_5980 & mul_34_17_n_6069)));
 assign mul_34_17_n_7105 = ((mul_34_17_n_5578 & mul_34_17_n_5746) | ((mul_34_17_n_5578 & mul_34_17_n_4248)
    | (mul_34_17_n_4248 & mul_34_17_n_5746)));
 assign mul_34_17_n_7104 = (mul_34_17_n_62 ^ mul_34_17_n_6666);
 assign mul_34_17_n_7103 = ((mul_34_17_n_5598 & mul_34_17_n_5732) | ((mul_34_17_n_5598 & mul_34_17_n_3060)
    | (mul_34_17_n_3060 & mul_34_17_n_5732)));
 assign mul_34_17_n_7101 = ((mul_34_17_n_5516 & mul_34_17_n_6044) | ((mul_34_17_n_5516 & mul_34_17_n_5913)
    | (mul_34_17_n_5913 & mul_34_17_n_6044)));
 assign mul_34_17_n_7100 = ((mul_34_17_n_5623 & mul_34_17_n_5743) | ((mul_34_17_n_5623 & mul_34_17_n_5622)
    | (mul_34_17_n_5622 & mul_34_17_n_5743)));
 assign mul_34_17_n_7099 = ((mul_34_17_n_5575 & mul_34_17_n_5728) | ((mul_34_17_n_5575 & mul_34_17_n_5576)
    | (mul_34_17_n_5576 & mul_34_17_n_5728)));
 assign mul_34_17_n_7098 = ((mul_34_17_n_5936 & mul_34_17_n_6050) | ((mul_34_17_n_5936 & mul_34_17_n_5939)
    | (mul_34_17_n_5939 & mul_34_17_n_6050)));
 assign mul_34_17_n_7097 = ((mul_34_17_n_4906 & mul_34_17_n_6140) | ((mul_34_17_n_4906 & mul_34_17_n_43)
    | (mul_34_17_n_43 & mul_34_17_n_6140)));
 assign mul_34_17_n_7095 = ((mul_34_17_n_5893 & mul_34_17_n_6071) | ((mul_34_17_n_5893 & mul_34_17_n_5985)
    | (mul_34_17_n_5985 & mul_34_17_n_6071)));
 assign mul_34_17_n_7094 = ~(mul_34_17_n_5156 ^ (mul_34_17_n_3800 ^ (mul_34_17_n_5157 ^ mul_34_17_n_3763)));
 assign mul_34_17_n_7093 = (mul_34_17_n_6373 ^ mul_34_17_n_6290);
 assign mul_34_17_n_7092 = ((mul_34_17_n_5918 & mul_34_17_n_6102) | ((mul_34_17_n_5918 & mul_34_17_n_5901)
    | (mul_34_17_n_5901 & mul_34_17_n_6102)));
 assign mul_34_17_n_7091 = ((mul_34_17_n_32 & mul_34_17_n_6203) | ((mul_34_17_n_32 & mul_34_17_n_5565)
    | (mul_34_17_n_5565 & mul_34_17_n_6203)));
 assign mul_34_17_n_7090 = ((mul_34_17_n_5961 & mul_34_17_n_6108) | ((mul_34_17_n_5961 & mul_34_17_n_6034)
    | (mul_34_17_n_6034 & mul_34_17_n_6108)));
 assign mul_34_17_n_7089 = ~(mul_34_17_n_5180 ^ (mul_34_17_n_4590 ^ (mul_34_17_n_5494 ^ mul_34_17_n_3695)));
 assign mul_34_17_n_7088 = ~(mul_34_17_n_5145 ^ (mul_34_17_n_3880 ^ (mul_34_17_n_5144 ^ mul_34_17_n_2813)));
 assign mul_34_17_n_7087 = ((mul_34_17_n_5556 & mul_34_17_n_5723) | ((mul_34_17_n_5556 & mul_34_17_n_5557)
    | (mul_34_17_n_5557 & mul_34_17_n_5723)));
 assign mul_34_17_n_7086 = (mul_34_17_n_6234 ^ mul_34_17_n_5705);
 assign mul_34_17_n_7085 = ((mul_34_17_n_5993 & mul_34_17_n_6110) | ((mul_34_17_n_5993 & mul_34_17_n_5204)
    | (mul_34_17_n_5204 & mul_34_17_n_6110)));
 assign mul_34_17_n_7084 = ~(mul_34_17_n_6432 ^ mul_34_17_n_5115);
 assign mul_34_17_n_7082 = ((mul_34_17_n_5613 & mul_34_17_n_89) | ((mul_34_17_n_5613 & mul_34_17_n_5560)
    | (mul_34_17_n_5560 & mul_34_17_n_89)));
 assign mul_34_17_n_7081 = ~(mul_34_17_n_5155 ^ (mul_34_17_n_3910 ^ (mul_34_17_n_5198 ^ mul_34_17_n_3838)));
 assign mul_34_17_n_7080 = ((mul_34_17_n_5915 & mul_34_17_n_6067) | ((mul_34_17_n_5915 & mul_34_17_n_5914)
    | (mul_34_17_n_5914 & mul_34_17_n_6067)));
 assign mul_34_17_n_7079 = ((mul_34_17_n_5528 & mul_34_17_n_8) | (mul_34_17_n_6440 & mul_34_17_n_5772));
 assign mul_34_17_n_7078 = ((mul_34_17_n_5507 & mul_34_17_n_6051) | ((mul_34_17_n_5507 & mul_34_17_n_3970)
    | (mul_34_17_n_3970 & mul_34_17_n_6051)));
 assign mul_34_17_n_7077 = ((mul_34_17_n_5902 & mul_34_17_n_5779) | ((mul_34_17_n_5902 & mul_34_17_n_5909)
    | (mul_34_17_n_5909 & mul_34_17_n_5779)));
 assign mul_34_17_n_7076 = ((mul_34_17_n_5539 & mul_34_17_n_5730) | ((mul_34_17_n_5539 & mul_34_17_n_5686)
    | (mul_34_17_n_5686 & mul_34_17_n_5730)));
 assign mul_34_17_n_7075 = ((mul_34_17_n_5674 & mul_34_17_n_6047) | ((mul_34_17_n_5674 & mul_34_17_n_3053)
    | (mul_34_17_n_3053 & mul_34_17_n_6047)));
 assign mul_34_17_n_7074 = (mul_34_17_n_6229 ^ mul_34_17_n_6370);
 assign mul_34_17_n_7073 = ((mul_34_17_n_5562 & mul_34_17_n_5726) | ((mul_34_17_n_5562 & mul_34_17_n_5563)
    | (mul_34_17_n_5563 & mul_34_17_n_5726)));
 assign mul_34_17_n_7072 = ((mul_34_17_n_5940 & mul_34_17_n_5739) | ((mul_34_17_n_5940 & mul_34_17_n_3031)
    | (mul_34_17_n_3031 & mul_34_17_n_5739)));
 assign mul_34_17_n_7071 = ((mul_34_17_n_5523 & mul_34_17_n_5439) | ((mul_34_17_n_5523 & mul_34_17_n_5524)
    | (mul_34_17_n_5524 & mul_34_17_n_5439)));
 assign mul_34_17_n_7070 = ((mul_34_17_n_5577 & mul_34_17_n_5442) | ((mul_34_17_n_5577 & mul_34_17_n_3491)
    | (mul_34_17_n_3491 & mul_34_17_n_5442)));
 assign mul_34_17_n_7069 = ((mul_34_17_n_140 & mul_34_17_n_5785) | ((mul_34_17_n_140 & mul_34_17_n_6008)
    | (mul_34_17_n_6008 & mul_34_17_n_5785)));
 assign mul_34_17_n_7068 = ((mul_34_17_n_127 & mul_34_17_n_5736) | ((mul_34_17_n_127 & mul_34_17_n_5604)
    | (mul_34_17_n_5604 & mul_34_17_n_5736)));
 assign mul_34_17_n_7067 = ~(mul_34_17_n_5192 ^ (mul_34_17_n_4691 ^ (mul_34_17_n_5191 ^ mul_34_17_n_4700)));
 assign mul_34_17_n_7066 = ((mul_34_17_n_5872 & mul_34_17_n_3979) | ((mul_34_17_n_5872 & mul_34_17_n_390)
    | (mul_34_17_n_390 & mul_34_17_n_3979)));
 assign mul_34_17_n_7065 = ((mul_34_17_n_5547 & mul_34_17_n_5441) | ((mul_34_17_n_5547 & mul_34_17_n_5548)
    | (mul_34_17_n_5548 & mul_34_17_n_5441)));
 assign mul_34_17_n_7064 = ((mul_34_17_n_5511 & mul_34_17_n_6073) | ((mul_34_17_n_5511 & mul_34_17_n_5991)
    | (mul_34_17_n_5991 & mul_34_17_n_6073)));
 assign mul_34_17_n_7062 = ~(mul_34_17_n_6430 ^ mul_34_17_n_5797);
 assign mul_34_17_n_7061 = ((mul_34_17_n_6021 & mul_34_17_n_5790) | ((mul_34_17_n_6021 & mul_34_17_n_3975)
    | (mul_34_17_n_3975 & mul_34_17_n_5790)));
 assign mul_34_17_n_7059 = ((mul_34_17_n_5620 & mul_34_17_n_6064) | ((mul_34_17_n_5620 & mul_34_17_n_5974)
    | (mul_34_17_n_5974 & mul_34_17_n_6064)));
 assign mul_34_17_n_7058 = ((mul_34_17_n_5958 & mul_34_17_n_6054) | ((mul_34_17_n_5958 & mul_34_17_n_5951)
    | (mul_34_17_n_5951 & mul_34_17_n_6054)));
 assign mul_34_17_n_7057 = ((mul_34_17_n_5591 & mul_34_17_n_5758) | ((mul_34_17_n_5591 & mul_34_17_n_5703)
    | (mul_34_17_n_5703 & mul_34_17_n_5758)));
 assign mul_34_17_n_7056 = ((mul_34_17_n_5573 & mul_34_17_n_5727) | ((mul_34_17_n_5573 & mul_34_17_n_4282)
    | (mul_34_17_n_4282 & mul_34_17_n_5727)));
 assign mul_34_17_n_7055 = ((mul_34_17_n_5986 & mul_34_17_n_6070) | ((mul_34_17_n_5986 & mul_34_17_n_5896)
    | (mul_34_17_n_5896 & mul_34_17_n_6070)));
 assign mul_34_17_n_7052 = ((mul_34_17_n_5585 & mul_34_17_n_6065) | ((mul_34_17_n_5585 & mul_34_17_n_5569)
    | (mul_34_17_n_5569 & mul_34_17_n_6065)));
 assign mul_34_17_n_7051 = ((mul_34_17_n_5581 & mul_34_17_n_5729) | ((mul_34_17_n_5581 & mul_34_17_n_5583)
    | (mul_34_17_n_5583 & mul_34_17_n_5729)));
 assign mul_34_17_n_7050 = ((mul_34_17_n_5935 & mul_34_17_n_6081) | ((mul_34_17_n_5935 & mul_34_17_n_46)
    | (mul_34_17_n_46 & mul_34_17_n_6081)));
 assign mul_34_17_n_7049 = ((mul_34_17_n_5550 & mul_34_17_n_5794) | ((mul_34_17_n_5550 & mul_34_17_n_5549)
    | (mul_34_17_n_5549 & mul_34_17_n_5794)));
 assign mul_34_17_n_6927 = ~mul_34_17_n_6926;
 assign mul_34_17_n_6924 = ~mul_34_17_n_190;
 assign mul_34_17_n_6903 = ~mul_34_17_n_6902;
 assign mul_34_17_n_6891 = ~(mul_34_17_n_6015 ^ mul_34_17_n_6016);
 assign mul_34_17_n_6890 = ~(mul_34_17_n_5931 ^ mul_34_17_n_5933);
 assign mul_34_17_n_6888 = ((mul_34_17_n_3958 | mul_34_17_n_2992) & (mul_34_17_n_6115 | mul_34_17_n_2867));
 assign mul_34_17_n_6887 = ~(mul_34_17_n_6487 & mul_34_17_n_6572);
 assign mul_34_17_n_6886 = ~(mul_34_17_n_6305 | mul_34_17_n_6675);
 assign mul_34_17_n_6885 = ~(mul_34_17_n_6561 & mul_34_17_n_136);
 assign mul_34_17_n_6884 = (mul_34_17_n_5558 ^ mul_34_17_n_5942);
 assign mul_34_17_n_6883 = ~(mul_34_17_n_5928 ^ mul_34_17_n_5938);
 assign mul_34_17_n_6882 = ~(mul_34_17_n_6307 | mul_34_17_n_5987);
 assign mul_34_17_n_6935 = ~(mul_34_17_n_6155 & mul_34_17_n_6356);
 assign mul_34_17_n_6876 = ~(mul_34_17_n_6304 | mul_34_17_n_6676);
 assign mul_34_17_n_6875 = ~(mul_34_17_n_6115 ^ mul_34_17_n_2867);
 assign mul_34_17_n_6934 = (mul_34_17_n_5888 ^ mul_34_17_n_4896);
 assign mul_34_17_n_6872 = ~(mul_34_17_n_6437 & mul_34_17_n_6364);
 assign mul_34_17_n_6871 = (mul_34_17_n_5938 ^ mul_34_17_n_5928);
 assign mul_34_17_n_6870 = (mul_34_17_n_5942 ^ mul_34_17_n_5558);
 assign mul_34_17_n_6867 = ~(mul_34_17_n_6016 ^ mul_34_17_n_6015);
 assign mul_34_17_n_6933 = ~(mul_34_17_n_6308 | mul_34_17_n_5108);
 assign mul_34_17_n_6864 = ~(mul_34_17_n_5932 ^ mul_34_17_n_5930);
 assign mul_34_17_n_6862 = (mul_34_17_n_5919 ^ mul_34_17_n_6097);
 assign mul_34_17_n_6861 = (mul_34_17_n_6032 ^ mul_34_17_n_5941);
 assign mul_34_17_n_6932 = (mul_34_17_n_5651 ^ mul_34_17_n_5753);
 assign mul_34_17_n_6860 = (mul_34_17_n_5756 ^ mul_34_17_n_5117);
 assign mul_34_17_n_6859 = (mul_34_17_n_5986 ^ mul_34_17_n_6070);
 assign mul_34_17_n_6858 = (mul_34_17_n_5761 ^ mul_34_17_n_5670);
 assign mul_34_17_n_6857 = (mul_34_17_n_5994 ^ mul_34_17_n_5996);
 assign mul_34_17_n_6856 = ~(mul_34_17_n_6076 ^ mul_34_17_n_4898);
 assign mul_34_17_n_6855 = (mul_34_17_n_5567 ^ mul_34_17_n_5675);
 assign mul_34_17_n_6854 = ~(mul_34_17_n_6119 & (mul_34_17_n_5840 & (mul_34_17_n_5864 & mul_34_17_n_6120)));
 assign mul_34_17_n_6853 = (mul_34_17_n_6009 ^ mul_34_17_n_6084);
 assign mul_34_17_n_6931 = ((mul_34_17_n_6116 & mul_34_17_n_3927) | (mul_34_17_n_6117 & mul_34_17_n_4844));
 assign mul_34_17_n_6852 = (mul_34_17_n_6017 ^ mul_34_17_n_6086);
 assign mul_34_17_n_6851 = (mul_34_17_n_6085 ^ mul_34_17_n_6014);
 assign mul_34_17_n_6850 = (mul_34_17_n_6090 ^ mul_34_17_n_6022);
 assign mul_34_17_n_6930 = (mul_34_17_n_6026 ^ mul_34_17_n_6094);
 assign mul_34_17_n_6929 = (mul_34_17_n_5429 ^ mul_34_17_n_6095);
 assign mul_34_17_n_6849 = (mul_34_17_n_5793 ^ mul_34_17_n_5621);
 assign mul_34_17_n_6928 = (mul_34_17_n_5572 ^ mul_34_17_n_5781);
 assign mul_34_17_n_6926 = ~(mul_34_17_n_5880 ^ mul_34_17_n_5417);
 assign mul_34_17_n_6848 = (mul_34_17_n_5805 ^ mul_34_17_n_5804);
 assign mul_34_17_n_6847 = (mul_34_17_n_6040 ^ mul_34_17_n_6027);
 assign mul_34_17_n_6846 = (mul_34_17_n_5766 ^ mul_34_17_n_5691);
 assign mul_34_17_n_6845 = (mul_34_17_n_6021 ^ mul_34_17_n_3975);
 assign mul_34_17_n_6844 = (mul_34_17_n_5636 ^ mul_34_17_n_5637);
 assign mul_34_17_n_6843 = (mul_34_17_n_5787 ^ mul_34_17_n_5618);
 assign mul_34_17_n_6842 = (mul_34_17_n_5693 ^ mul_34_17_n_5765);
 assign mul_34_17_n_6841 = (mul_34_17_n_6004 ^ mul_34_17_n_6112);
 assign mul_34_17_n_6840 = (mul_34_17_n_5910 ^ mul_34_17_n_5960);
 assign mul_34_17_n_6839 = ~(mul_34_17_n_5807 ^ mul_34_17_n_5502);
 assign mul_34_17_n_6838 = (mul_34_17_n_5976 ^ mul_34_17_n_5978);
 assign mul_34_17_n_6837 = ~(mul_34_17_n_5903 ^ mul_34_17_n_5894);
 assign mul_34_17_n_6836 = (mul_34_17_n_5971 ^ mul_34_17_n_5975);
 assign mul_34_17_n_6835 = (mul_34_17_n_3024 ^ mul_34_17_n_6038);
 assign mul_34_17_n_6834 = ~(mul_34_17_n_6104 ^ mul_34_17_n_4893);
 assign mul_34_17_n_6832 = ~(mul_34_17_n_6183 | mul_34_17_n_6178);
 assign mul_34_17_n_6925 = (mul_34_17_n_5984 ^ mul_34_17_n_5892);
 assign mul_34_17_n_6831 = (mul_34_17_n_5955 ^ mul_34_17_n_6103);
 assign mul_34_17_n_6830 = ~(mul_34_17_n_6078 ^ mul_34_17_n_3033);
 assign mul_34_17_n_6829 = (mul_34_17_n_140 ^ mul_34_17_n_6008);
 assign mul_34_17_n_6828 = (mul_34_17_n_137 ^ mul_34_17_n_6005);
 assign mul_34_17_n_6827 = (mul_34_17_n_5616 ^ mul_34_17_n_5786);
 assign mul_34_17_n_6826 = ~(mul_34_17_n_6402 & mul_34_17_n_6682);
 assign mul_34_17_n_6825 = (mul_34_17_n_5545 ^ mul_34_17_n_5543);
 assign mul_34_17_n_6824 = (mul_34_17_n_6012 ^ mul_34_17_n_5998);
 assign mul_34_17_n_6823 = (mul_34_17_n_5740 ^ mul_34_17_n_5692);
 assign mul_34_17_n_6822 = (mul_34_17_n_129 ^ mul_34_17_n_131);
 assign mul_34_17_n_6821 = (mul_34_17_n_5660 ^ mul_34_17_n_5601);
 assign mul_34_17_n_6820 = (mul_34_17_n_5959 ^ mul_34_17_n_5956);
 assign mul_34_17_n_6819 = (mul_34_17_n_6106 ^ mul_34_17_n_6006);
 assign mul_34_17_n_6818 = (mul_34_17_n_5652 ^ mul_34_17_n_5449);
 assign mul_34_17_n_6817 = (mul_34_17_n_4391 ^ mul_34_17_n_6052);
 assign mul_34_17_n_6816 = (mul_34_17_n_5701 ^ mul_34_17_n_5700);
 assign mul_34_17_n_6923 = ((mul_34_17_n_3055 & mul_34_17_n_6059) | ((mul_34_17_n_3055 & mul_34_17_n_3943)
    | (mul_34_17_n_3943 & mul_34_17_n_6059)));
 assign mul_34_17_n_6922 = ((mul_34_17_n_3172 & mul_34_17_n_5881) | ((mul_34_17_n_3172 & mul_34_17_n_3634)
    | (mul_34_17_n_3634 & mul_34_17_n_5881)));
 assign mul_34_17_n_6815 = ~(mul_34_17_n_6408 | mul_34_17_n_6687);
 assign mul_34_17_n_6921 = ~(mul_34_17_n_6408 & mul_34_17_n_6687);
 assign mul_34_17_n_6814 = ~(mul_34_17_n_6403 & mul_34_17_n_5465);
 assign mul_34_17_n_6920 = ((mul_34_17_n_5499 & mul_34_17_n_5797) | ((mul_34_17_n_5499 & mul_34_17_n_4825)
    | (mul_34_17_n_4825 & mul_34_17_n_5797)));
 assign mul_34_17_n_6919 = ((mul_34_17_n_3964 & mul_34_17_n_6082) | ((mul_34_17_n_3964 & mul_34_17_n_4840)
    | (mul_34_17_n_4840 & mul_34_17_n_6082)));
 assign mul_34_17_n_6918 = ((mul_34_17_n_5503 & mul_34_17_n_5451) | (mul_34_17_n_5833 & mul_34_17_n_5403));
 assign mul_34_17_n_6917 = ((mul_34_17_n_4888 & mul_34_17_n_5784) | ((mul_34_17_n_4888 & mul_34_17_n_4178)
    | (mul_34_17_n_4178 & mul_34_17_n_5784)));
 assign mul_34_17_n_6916 = ((mul_34_17_n_4891 & mul_34_17_n_5800) | ((mul_34_17_n_4891 & mul_34_17_n_4442)
    | (mul_34_17_n_4442 & mul_34_17_n_5800)));
 assign mul_34_17_n_6915 = ~(mul_34_17_n_6082 ^ mul_34_17_n_5339);
 assign mul_34_17_n_6914 = ((mul_34_17_n_4897 & mul_34_17_n_6089) | ((mul_34_17_n_4897 & mul_34_17_n_3512)
    | (mul_34_17_n_3512 & mul_34_17_n_6089)));
 assign mul_34_17_n_6913 = ((mul_34_17_n_4902 & mul_34_17_n_5755) | ((mul_34_17_n_4902 & mul_34_17_n_3930)
    | (mul_34_17_n_3930 & mul_34_17_n_5755)));
 assign mul_34_17_n_6912 = (mul_34_17_n_5780 ^ mul_34_17_n_3961);
 assign mul_34_17_n_6911 = ((mul_34_17_n_4836 & mul_34_17_n_6092) | ((mul_34_17_n_4836 & mul_34_17_n_3037)
    | (mul_34_17_n_3037 & mul_34_17_n_6092)));
 assign mul_34_17_n_6910 = (mul_34_17_n_5775 ^ mul_34_17_n_5536);
 assign mul_34_17_n_6909 = ((mul_34_17_n_5420 & mul_34_17_n_6100) | ((mul_34_17_n_5420 & mul_34_17_n_4436)
    | (mul_34_17_n_4436 & mul_34_17_n_6100)));
 assign mul_34_17_n_6908 = ((mul_34_17_n_3940 & mul_34_17_n_3040) | (mul_34_17_n_5819 & mul_34_17_n_4876));
 assign mul_34_17_n_6907 = (mul_34_17_n_6072 ^ mul_34_17_n_5990);
 assign mul_34_17_n_6906 = ((mul_34_17_n_3970 & mul_34_17_n_125) | ((mul_34_17_n_3970 & mul_34_17_n_4842)
    | (mul_34_17_n_4842 & mul_34_17_n_125)));
 assign mul_34_17_n_6905 = ((mul_34_17_n_4901 & mul_34_17_n_5877) | ((mul_34_17_n_4901 & mul_34_17_n_4831)
    | (mul_34_17_n_4831 & mul_34_17_n_5877)));
 assign mul_34_17_n_6904 = ((mul_34_17_n_4827 & mul_34_17_n_5880) | ((mul_34_17_n_4827 & mul_34_17_n_3041)
    | (mul_34_17_n_3041 & mul_34_17_n_5880)));
 assign mul_34_17_n_6902 = ~((mul_34_17_n_3975 | mul_34_17_n_3932) & (mul_34_17_n_5878 | mul_34_17_n_67));
 assign mul_34_17_n_6901 = ((mul_34_17_n_3931 & mul_34_17_n_6114) | ((mul_34_17_n_3931 & mul_34_17_n_3058)
    | (mul_34_17_n_3058 & mul_34_17_n_6114)));
 assign mul_34_17_n_6900 = ~((mul_34_17_n_3060 & mul_34_17_n_3942) | (mul_34_17_n_5883 & mul_34_17_n_4880));
 assign mul_34_17_n_6899 = (mul_34_17_n_6098 ^ mul_34_17_n_103);
 assign mul_34_17_n_6898 = (mul_34_17_n_5764 ^ mul_34_17_n_5689);
 assign mul_34_17_n_6897 = ((mul_34_17_n_5111 & mul_34_17_n_5721) | ((mul_34_17_n_5111 & mul_34_17_n_4372)
    | (mul_34_17_n_4372 & mul_34_17_n_5721)));
 assign mul_34_17_n_6896 = ((mul_34_17_n_3500 & mul_34_17_n_6039) | ((mul_34_17_n_3500 & mul_34_17_n_3027)
    | (mul_34_17_n_3027 & mul_34_17_n_6039)));
 assign mul_34_17_n_6895 = ~(mul_34_17_n_6089 ^ mul_34_17_n_5812);
 assign mul_34_17_n_6894 = ~(mul_34_17_n_6091 ^ mul_34_17_n_5332);
 assign mul_34_17_n_6893 = ~(mul_34_17_n_5394 ^ mul_34_17_n_6113);
 assign mul_34_17_n_6813 = ~mul_34_17_n_6812;
 assign mul_34_17_n_6801 = ~mul_34_17_n_6800;
 assign mul_34_17_n_6791 = ~mul_34_17_n_6792;
 assign mul_34_17_n_6784 = ~mul_34_17_n_6783;
 assign mul_34_17_n_6782 = ~mul_34_17_n_6781;
 assign mul_34_17_n_6767 = ~(mul_34_17_n_5505 ^ mul_34_17_n_5886);
 assign mul_34_17_n_6812 = ~(mul_34_17_n_5888 ^ mul_34_17_n_4896);
 assign mul_34_17_n_6764 = ~(mul_34_17_n_6088 ^ mul_34_17_n_5528);
 assign mul_34_17_n_6763 = (mul_34_17_n_6062 ^ mul_34_17_n_5969);
 assign mul_34_17_n_6762 = (mul_34_17_n_5610 ^ mul_34_17_n_5738);
 assign mul_34_17_n_6761 = (mul_34_17_n_6043 ^ mul_34_17_n_6024);
 assign mul_34_17_n_6811 = (mul_34_17_n_5727 ^ mul_34_17_n_4282);
 assign mul_34_17_n_6760 = (mul_34_17_n_6045 ^ mul_34_17_n_5907);
 assign mul_34_17_n_6810 = (mul_34_17_n_5729 ^ mul_34_17_n_5583);
 assign mul_34_17_n_6759 = (mul_34_17_n_5799 ^ mul_34_17_n_5537);
 assign mul_34_17_n_6758 = (mul_34_17_n_5918 ^ mul_34_17_n_5901);
 assign mul_34_17_n_6809 = (mul_34_17_n_5974 ^ mul_34_17_n_6064);
 assign mul_34_17_n_6757 = (mul_34_17_n_6060 ^ mul_34_17_n_3023);
 assign mul_34_17_n_6756 = (mul_34_17_n_5760 ^ mul_34_17_n_5541);
 assign mul_34_17_n_6755 = (mul_34_17_n_5954 ^ mul_34_17_n_6055);
 assign mul_34_17_n_6754 = (mul_34_17_n_5951 ^ mul_34_17_n_6054);
 assign mul_34_17_n_6753 = (mul_34_17_n_5742 ^ mul_34_17_n_3962);
 assign mul_34_17_n_6752 = (mul_34_17_n_5622 ^ mul_34_17_n_5743);
 assign mul_34_17_n_6751 = (mul_34_17_n_56 ^ mul_34_17_n_5609);
 assign mul_34_17_n_6750 = (mul_34_17_n_5628 ^ mul_34_17_n_105);
 assign mul_34_17_n_6749 = (mul_34_17_n_5653 ^ mul_34_17_n_5716);
 assign mul_34_17_n_6748 = (mul_34_17_n_5523 ^ mul_34_17_n_5439);
 assign mul_34_17_n_6747 = (mul_34_17_n_75 ^ mul_34_17_n_6053);
 assign mul_34_17_n_6808 = ~(mul_34_17_n_5125 ^ mul_34_17_n_5881);
 assign mul_34_17_n_6746 = (mul_34_17_n_6099 ^ mul_34_17_n_5929);
 assign mul_34_17_n_6745 = (mul_34_17_n_5711 ^ mul_34_17_n_5773);
 assign mul_34_17_n_6744 = (mul_34_17_n_6018 ^ mul_34_17_n_6011);
 assign mul_34_17_n_6743 = (mul_34_17_n_5940 ^ mul_34_17_n_3031);
 assign mul_34_17_n_6742 = (mul_34_17_n_5626 ^ mul_34_17_n_5745);
 assign mul_34_17_n_6741 = (mul_34_17_n_5709 ^ mul_34_17_n_5770);
 assign mul_34_17_n_6740 = (mul_34_17_n_5774 ^ mul_34_17_n_5555);
 assign mul_34_17_n_6739 = (mul_34_17_n_5924 ^ mul_34_17_n_5925);
 assign mul_34_17_n_6738 = (mul_34_17_n_5908 ^ mul_34_17_n_6049);
 assign mul_34_17_n_6737 = (mul_34_17_n_5939 ^ mul_34_17_n_5936);
 assign mul_34_17_n_6736 = (mul_34_17_n_127 ^ mul_34_17_n_5736);
 assign mul_34_17_n_6735 = (mul_34_17_n_5754 ^ mul_34_17_n_5639);
 assign mul_34_17_n_6734 = (mul_34_17_n_5735 ^ mul_34_17_n_5600);
 assign mul_34_17_n_6733 = ~(mul_34_17_n_6046 ^ mul_34_17_n_3053);
 assign mul_34_17_n_6807 = ~(mul_34_17_n_5989 ^ mul_34_17_n_5416);
 assign mul_34_17_n_6732 = (mul_34_17_n_5962 ^ mul_34_17_n_6058);
 assign mul_34_17_n_6731 = (mul_34_17_n_5646 ^ mul_34_17_n_5751);
 assign mul_34_17_n_6730 = ~(mul_34_17_n_6096 ^ mul_34_17_n_5642);
 assign mul_34_17_n_6729 = (mul_34_17_n_5612 ^ mul_34_17_n_5559);
 assign mul_34_17_n_6728 = ~(mul_34_17_n_5915 ^ mul_34_17_n_5914);
 assign mul_34_17_n_6727 = (mul_34_17_n_5748 ^ mul_34_17_n_5634);
 assign mul_34_17_n_6726 = (mul_34_17_n_5663 ^ mul_34_17_n_5759);
 assign mul_34_17_n_6725 = (mul_34_17_n_5686 ^ mul_34_17_n_5730);
 assign mul_34_17_n_6724 = (mul_34_17_n_49 ^ mul_34_17_n_113);
 assign mul_34_17_n_6723 = (mul_34_17_n_5979 ^ mul_34_17_n_6068);
 assign mul_34_17_n_6806 = (mul_34_17_n_5569 ^ mul_34_17_n_6065);
 assign mul_34_17_n_6805 = (mul_34_17_n_5717 ^ mul_34_17_n_5662);
 assign mul_34_17_n_6722 = (mul_34_17_n_5676 ^ mul_34_17_n_5762);
 assign mul_34_17_n_6721 = (mul_34_17_n_5592 ^ mul_34_17_n_5594);
 assign mul_34_17_n_6720 = (mul_34_17_n_5643 ^ mul_34_17_n_5750);
 assign mul_34_17_n_6719 = (mul_34_17_n_6063 ^ mul_34_17_n_5972);
 assign mul_34_17_n_6718 = (mul_34_17_n_5752 ^ mul_34_17_n_4887);
 assign mul_34_17_n_6717 = (mul_34_17_n_5801 ^ mul_34_17_n_5526);
 assign mul_34_17_n_6716 = (mul_34_17_n_5796 ^ mul_34_17_n_5659);
 assign mul_34_17_n_6715 = (mul_34_17_n_5521 ^ mul_34_17_n_5681);
 assign mul_34_17_n_6714 = (mul_34_17_n_4412 ^ mul_34_17_n_6048);
 assign mul_34_17_n_6713 = (mul_34_17_n_5614 ^ mul_34_17_n_5889);
 assign mul_34_17_n_6712 = (mul_34_17_n_5724 ^ mul_34_17_n_5566);
 assign mul_34_17_n_6711 = (mul_34_17_n_6042 ^ mul_34_17_n_4895);
 assign mul_34_17_n_6710 = (mul_34_17_n_5737 ^ mul_34_17_n_5109);
 assign mul_34_17_n_6709 = (mul_34_17_n_6083 ^ mul_34_17_n_5899);
 assign mul_34_17_n_6708 = (mul_34_17_n_6080 ^ mul_34_17_n_6007);
 assign mul_34_17_n_6707 = (mul_34_17_n_5945 ^ mul_34_17_n_5887);
 assign mul_34_17_n_6706 = (mul_34_17_n_5965 ^ mul_34_17_n_5981);
 assign mul_34_17_n_6705 = (mul_34_17_n_5935 ^ mul_34_17_n_46);
 assign mul_34_17_n_6804 = (mul_34_17_n_5948 ^ mul_34_17_n_6057);
 assign mul_34_17_n_6704 = (mul_34_17_n_5631 ^ mul_34_17_n_5771);
 assign mul_34_17_n_6703 = (mul_34_17_n_6087 ^ mul_34_17_n_4892);
 assign mul_34_17_n_6702 = (mul_34_17_n_5571 ^ mul_34_17_n_5795);
 assign mul_34_17_n_6701 = (mul_34_17_n_5728 ^ mul_34_17_n_5576);
 assign mul_34_17_n_6700 = (mul_34_17_n_5562 ^ mul_34_17_n_5726);
 assign mul_34_17_n_6699 = (mul_34_17_n_5702 ^ mul_34_17_n_5590);
 assign mul_34_17_n_6698 = (mul_34_17_n_5598 ^ mul_34_17_n_3060);
 assign mul_34_17_n_6697 = (mul_34_17_n_6108 ^ mul_34_17_n_5961);
 assign mul_34_17_n_6696 = (mul_34_17_n_5540 ^ mul_34_17_n_5114);
 assign mul_34_17_n_6695 = (mul_34_17_n_5721 ^ mul_34_17_n_4372);
 assign mul_34_17_n_6694 = (mul_34_17_n_5549 ^ mul_34_17_n_5794);
 assign mul_34_17_n_6693 = (mul_34_17_n_5909 ^ mul_34_17_n_5902);
 assign mul_34_17_n_6803 = (mul_34_17_n_5722 ^ mul_34_17_n_5553);
 assign mul_34_17_n_6692 = (mul_34_17_n_5746 ^ mul_34_17_n_4248);
 assign mul_34_17_n_6691 = (mul_34_17_n_5548 ^ mul_34_17_n_5441);
 assign mul_34_17_n_6690 = (mul_34_17_n_5720 ^ mul_34_17_n_5542);
 assign mul_34_17_n_6689 = (mul_34_17_n_5723 ^ mul_34_17_n_5557);
 assign mul_34_17_n_6802 = ~(mul_34_17_n_5800 ^ mul_34_17_n_5501);
 assign mul_34_17_n_6800 = ~(mul_34_17_n_5811 ^ mul_34_17_n_3523);
 assign mul_34_17_n_6798 = ~(mul_34_17_n_6059 ^ mul_34_17_n_5330);
 assign mul_34_17_n_6797 = ((mul_34_17_n_5115 & mul_34_17_n_5446) | ((mul_34_17_n_5115 & mul_34_17_n_3380)
    | (mul_34_17_n_3380 & mul_34_17_n_5446)));
 assign mul_34_17_n_6796 = (mul_34_17_n_5916 ^ mul_34_17_n_6056);
 assign mul_34_17_n_6795 = (mul_34_17_n_6044 ^ mul_34_17_n_5913);
 assign mul_34_17_n_6794 = ~(mul_34_17_n_125 ^ mul_34_17_n_5389);
 assign mul_34_17_n_6793 = (mul_34_17_n_5565 ^ mul_34_17_n_32);
 assign mul_34_17_n_6792 = (mul_34_17_n_3970 ^ mul_34_17_n_6051);
 assign mul_34_17_n_6790 = (mul_34_17_n_5625 ^ mul_34_17_n_5744);
 assign mul_34_17_n_6789 = ~(mul_34_17_n_5755 ^ mul_34_17_n_5813);
 assign mul_34_17_n_6788 = (mul_34_17_n_5629 ^ mul_34_17_n_5627);
 assign mul_34_17_n_6787 = ((mul_34_17_n_4220 & mul_34_17_n_5734) | ((mul_34_17_n_4220 & mul_34_17_n_4350)
    | (mul_34_17_n_4350 & mul_34_17_n_5734)));
 assign mul_34_17_n_6786 = ~(mul_34_17_n_5096 ^ mul_34_17_n_5733);
 assign mul_34_17_n_6785 = (mul_34_17_n_5747 ^ mul_34_17_n_5635);
 assign mul_34_17_n_6783 = ((mul_34_17_n_5113 & mul_34_17_n_4668) | ((mul_34_17_n_5113 & mul_34_17_n_3364)
    | (mul_34_17_n_3364 & mul_34_17_n_4668)));
 assign mul_34_17_n_6781 = ((mul_34_17_n_5108 & mul_34_17_n_5445) | ((mul_34_17_n_5108 & mul_34_17_n_2834)
    | (mul_34_17_n_2834 & mul_34_17_n_5445)));
 assign mul_34_17_n_6780 = ~(mul_34_17_n_6039 ^ mul_34_17_n_5021);
 assign mul_34_17_n_6779 = ~(mul_34_17_n_5809 ^ mul_34_17_n_5749);
 assign mul_34_17_n_6778 = ((mul_34_17_n_4890 & mul_34_17_n_5749) | ((mul_34_17_n_4890 & mul_34_17_n_3963)
    | (mul_34_17_n_3963 & mul_34_17_n_5749)));
 assign mul_34_17_n_6777 = ((mul_34_17_n_3054 & mul_34_17_n_6066) | ((mul_34_17_n_3054 & mul_34_17_n_4099)
    | (mul_34_17_n_4099 & mul_34_17_n_6066)));
 assign mul_34_17_n_6776 = ~(mul_34_17_n_5810 ^ mul_34_17_n_5784);
 assign mul_34_17_n_6686 = ~mul_34_17_n_6687;
 assign mul_34_17_n_6681 = ~mul_34_17_n_6680;
 assign mul_34_17_n_6679 = ~mul_34_17_n_6678;
 assign mul_34_17_n_6675 = ~mul_34_17_n_6676;
 assign mul_34_17_n_6662 = ~mul_34_17_n_71;
 assign mul_34_17_n_6661 = ~mul_34_17_n_6660;
 assign mul_34_17_n_6653 = ~mul_34_17_n_6652;
 assign mul_34_17_n_6647 = ~mul_34_17_n_6646;
 assign mul_34_17_n_6645 = ~mul_34_17_n_6644;
 assign mul_34_17_n_6643 = ~mul_34_17_n_6642;
 assign mul_34_17_n_6638 = ~mul_34_17_n_6637;
 assign mul_34_17_n_6635 = ~mul_34_17_n_6634;
 assign mul_34_17_n_6603 = ~mul_34_17_n_6604;
 assign mul_34_17_n_6598 = ~mul_34_17_n_6597;
 assign mul_34_17_n_6596 = ~mul_34_17_n_6595;
 assign mul_34_17_n_6573 = ~mul_34_17_n_6572;
 assign mul_34_17_n_6568 = ~mul_34_17_n_6567;
 assign mul_34_17_n_6562 = ~mul_34_17_n_6561;
 assign mul_34_17_n_6521 = ~mul_34_17_n_6522;
 assign mul_34_17_n_6519 = ~mul_34_17_n_6520;
 assign mul_34_17_n_6512 = ~mul_34_17_n_6513;
 assign mul_34_17_n_6493 = ~mul_34_17_n_136;
 assign mul_34_17_n_6491 = ~mul_34_17_n_6492;
 assign mul_34_17_n_6490 = ~mul_34_17_n_6489;
 assign mul_34_17_n_6486 = ~mul_34_17_n_6487;
 assign mul_34_17_n_6476 = ~mul_34_17_n_6477;
 assign mul_34_17_n_6456 = ~mul_34_17_n_6457;
 assign mul_34_17_n_6455 = ~mul_34_17_n_145;
 assign mul_34_17_n_6451 = ~(mul_34_17_n_5879 & mul_34_17_n_5414);
 assign mul_34_17_n_6450 = ~(mul_34_17_n_5879 | mul_34_17_n_5414);
 assign mul_34_17_n_6449 = ~(mul_34_17_n_5127 ^ mul_34_17_n_3071);
 assign mul_34_17_n_6448 = ~(mul_34_17_n_5883 & mul_34_17_n_5415);
 assign mul_34_17_n_6447 = ~(mul_34_17_n_5883 | mul_34_17_n_5415);
 assign mul_34_17_n_6446 = ~(mul_34_17_n_5641 & mul_34_17_n_6096);
 assign mul_34_17_n_6445 = ~(mul_34_17_n_5887 & mul_34_17_n_6010);
 assign mul_34_17_n_6444 = ~(mul_34_17_n_5880 & mul_34_17_n_5417);
 assign mul_34_17_n_6443 = ~(mul_34_17_n_5880 | mul_34_17_n_5417);
 assign mul_34_17_n_6442 = ~(mul_34_17_n_6117 & mul_34_17_n_4844);
 assign mul_34_17_n_6441 = ~(mul_34_17_n_5989 | mul_34_17_n_5416);
 assign mul_34_17_n_6440 = ~(mul_34_17_n_6088 & mul_34_17_n_5527);
 assign mul_34_17_n_6439 = ~(mul_34_17_n_5989 & mul_34_17_n_5416);
 assign mul_34_17_n_6438 = ~(mul_34_17_n_5135 & mul_34_17_n_5898);
 assign mul_34_17_n_6437 = ~(mul_34_17_n_5136 & mul_34_17_n_5897);
 assign mul_34_17_n_6436 = ~(mul_34_17_n_6116 & mul_34_17_n_3927);
 assign mul_34_17_n_6435 = ~(mul_34_17_n_5877 & mul_34_17_n_6025);
 assign mul_34_17_n_6434 = ~(mul_34_17_n_5877 | mul_34_17_n_6025);
 assign mul_34_17_n_6688 = ~(mul_34_17_n_5421 ^ mul_34_17_n_3972);
 assign mul_34_17_n_6687 = ((mul_34_17_n_4851 & mul_34_17_n_3927) | ((mul_34_17_n_4851 & mul_34_17_n_3087)
    | (mul_34_17_n_3087 & mul_34_17_n_3927)));
 assign mul_34_17_n_6433 = ~(mul_34_17_n_6000 & mul_34_17_n_6006);
 assign mul_34_17_n_6432 = (mul_34_17_n_5446 ^ mul_34_17_n_3380);
 assign mul_34_17_n_6685 = ~(mul_34_17_n_5438 ^ mul_34_17_n_3973);
 assign mul_34_17_n_6684 = ~(mul_34_17_n_5434 ^ mul_34_17_n_3075);
 assign mul_34_17_n_6683 = ~(mul_34_17_n_5430 ^ mul_34_17_n_3980);
 assign mul_34_17_n_6682 = ~(mul_34_17_n_5173 ^ mul_34_17_n_4872);
 assign mul_34_17_n_6680 = ~(mul_34_17_n_5431 ^ mul_34_17_n_2809);
 assign mul_34_17_n_6678 = ~(mul_34_17_n_5436 ^ mul_34_17_n_3067);
 assign mul_34_17_n_6431 = ~(mul_34_17_n_5965 & mul_34_17_n_5981);
 assign mul_34_17_n_6430 = ~(mul_34_17_n_5499 ^ mul_34_17_n_4825);
 assign mul_34_17_n_6677 = ~(mul_34_17_n_5326 ^ mul_34_17_n_4058);
 assign mul_34_17_n_6676 = ~(mul_34_17_n_5390 ^ mul_34_17_n_5);
 assign mul_34_17_n_6674 = ~(mul_34_17_n_5325 ^ mul_34_17_n_4031);
 assign mul_34_17_n_6429 = (mul_34_17_n_390 ^ mul_34_17_n_3979);
 assign mul_34_17_n_6428 = ~(mul_34_17_n_5949 & mul_34_17_n_5952);
 assign mul_34_17_n_6427 = (mul_34_17_n_4436 ^ mul_34_17_n_5420);
 assign mul_34_17_n_6673 = ((mul_34_17_n_5396 & mul_34_17_n_3960) | (mul_34_17_n_5408 & mul_34_17_n_4));
 assign mul_34_17_n_6426 = (mul_34_17_n_5457 ^ mul_34_17_n_4181);
 assign mul_34_17_n_6671 = ~(mul_34_17_n_5233 ^ mul_34_17_n_3405);
 assign mul_34_17_n_6425 = ~(mul_34_17_n_5494 ^ mul_34_17_n_3695);
 assign mul_34_17_n_6670 = ~(mul_34_17_n_5485 ^ mul_34_17_n_4747);
 assign mul_34_17_n_6668 = ~(mul_34_17_n_5236 ^ mul_34_17_n_3529);
 assign mul_34_17_n_6667 = ~(mul_34_17_n_5379 ^ mul_34_17_n_4787);
 assign mul_34_17_n_6666 = ~(mul_34_17_n_4866 ^ mul_34_17_n_5237);
 assign mul_34_17_n_6665 = ~(mul_34_17_n_5254 ^ mul_34_17_n_4299);
 assign mul_34_17_n_6664 = ~(mul_34_17_n_5260 ^ mul_34_17_n_4630);
 assign mul_34_17_n_6663 = ~(mul_34_17_n_4942 ^ mul_34_17_n_3728);
 assign mul_34_17_n_6660 = ~(mul_34_17_n_5377 ^ mul_34_17_n_4290);
 assign mul_34_17_n_6659 = ~(mul_34_17_n_5263 ^ mul_34_17_n_4855);
 assign mul_34_17_n_6657 = ~(mul_34_17_n_5293 ^ mul_34_17_n_5113);
 assign mul_34_17_n_6655 = ~(mul_34_17_n_5346 ^ mul_34_17_n_3058);
 assign mul_34_17_n_6654 = ~(mul_34_17_n_5432 ^ mul_34_17_n_3982);
 assign mul_34_17_n_6652 = ~(mul_34_17_n_5437 ^ mul_34_17_n_3978);
 assign mul_34_17_n_6650 = ~(mul_34_17_n_5262 ^ mul_34_17_n_4216);
 assign mul_34_17_n_6649 = ((mul_34_17_n_4850 & mul_34_17_n_5452) | ((mul_34_17_n_4850 & mul_34_17_n_3300)
    | (mul_34_17_n_3300 & mul_34_17_n_5452)));
 assign mul_34_17_n_6648 = ~(mul_34_17_n_5342 ^ mul_34_17_n_4761);
 assign mul_34_17_n_6646 = ~(mul_34_17_n_5418 ^ mul_34_17_n_3985);
 assign mul_34_17_n_6644 = ~(mul_34_17_n_5419 ^ mul_34_17_n_3966);
 assign mul_34_17_n_6424 = (mul_34_17_n_5490 ^ mul_34_17_n_4468);
 assign mul_34_17_n_6423 = (mul_34_17_n_5152 ^ mul_34_17_n_3716);
 assign mul_34_17_n_6642 = ~(mul_34_17_n_5110 ^ mul_34_17_n_3969);
 assign mul_34_17_n_6641 = ((mul_34_17_n_3476 & mul_34_17_n_5444) | ((mul_34_17_n_3476 & mul_34_17_n_3559)
    | (mul_34_17_n_3559 & mul_34_17_n_5444)));
 assign mul_34_17_n_6422 = (mul_34_17_n_5476 ^ mul_34_17_n_3532);
 assign mul_34_17_n_6421 = (mul_34_17_n_5489 ^ mul_34_17_n_4116);
 assign mul_34_17_n_6640 = ~(mul_34_17_n_5042 ^ mul_34_17_n_4173);
 assign mul_34_17_n_6639 = (mul_34_17_n_5470 ^ mul_34_17_n_4687);
 assign mul_34_17_n_6637 = ~(mul_34_17_n_5337 ^ mul_34_17_n_3036);
 assign mul_34_17_n_6636 = ~(mul_34_17_n_5426 ^ mul_34_17_n_3971);
 assign mul_34_17_n_6634 = ~(mul_34_17_n_5423 ^ mul_34_17_n_3072);
 assign mul_34_17_n_6633 = ~(mul_34_17_n_5060 ^ mul_34_17_n_3374);
 assign mul_34_17_n_6632 = ~(mul_34_17_n_5221 ^ mul_34_17_n_4201);
 assign mul_34_17_n_6631 = ~(mul_34_17_n_5422 ^ mul_34_17_n_3974);
 assign mul_34_17_n_6630 = ~(mul_34_17_n_5264 ^ mul_34_17_n_4648);
 assign mul_34_17_n_6420 = ~(mul_34_17_n_5177 ^ mul_34_17_n_4726);
 assign mul_34_17_n_6629 = ~(mul_34_17_n_5297 ^ mul_34_17_n_4867);
 assign mul_34_17_n_6628 = ~(mul_34_17_n_5387 ^ mul_34_17_n_3148);
 assign mul_34_17_n_6627 = ~(mul_34_17_n_5307 ^ mul_34_17_n_4131);
 assign mul_34_17_n_6626 = ~(mul_34_17_n_5311 ^ mul_34_17_n_4721);
 assign mul_34_17_n_6625 = (mul_34_17_n_5492 ^ mul_34_17_n_4429);
 assign mul_34_17_n_6624 = (mul_34_17_n_5466 ^ mul_34_17_n_3860);
 assign mul_34_17_n_6623 = ~(mul_34_17_n_5306 ^ mul_34_17_n_3305);
 assign mul_34_17_n_6622 = (mul_34_17_n_5463 ^ mul_34_17_n_3391);
 assign mul_34_17_n_6621 = (mul_34_17_n_5478 ^ mul_34_17_n_3115);
 assign mul_34_17_n_6620 = ~(mul_34_17_n_5341 ^ mul_34_17_n_4575);
 assign mul_34_17_n_6619 = ~(mul_34_17_n_5309 ^ mul_34_17_n_4742);
 assign mul_34_17_n_6618 = ~(mul_34_17_n_5083 ^ mul_34_17_n_3872);
 assign mul_34_17_n_6617 = ~(mul_34_17_n_5301 ^ mul_34_17_n_4718);
 assign mul_34_17_n_6616 = ~(mul_34_17_n_4937 ^ mul_34_17_n_3961);
 assign mul_34_17_n_6615 = ~(mul_34_17_n_5312 ^ mul_34_17_n_4772);
 assign mul_34_17_n_6614 = ~(mul_34_17_n_5040 ^ mul_34_17_n_4698);
 assign mul_34_17_n_6613 = ~(mul_34_17_n_5295 ^ mul_34_17_n_4871);
 assign mul_34_17_n_6611 = ~(mul_34_17_n_5048 ^ mul_34_17_n_4817);
 assign mul_34_17_n_6610 = ~(mul_34_17_n_5294 ^ mul_34_17_n_4694);
 assign mul_34_17_n_6419 = (mul_34_17_n_5469 ^ mul_34_17_n_4736);
 assign mul_34_17_n_6609 = ~(mul_34_17_n_5292 ^ mul_34_17_n_4719);
 assign mul_34_17_n_6608 = ~(mul_34_17_n_5380 ^ mul_34_17_n_4766);
 assign mul_34_17_n_6607 = ~(mul_34_17_n_5265 ^ mul_34_17_n_4470);
 assign mul_34_17_n_6606 = ~(mul_34_17_n_5322 ^ mul_34_17_n_4345);
 assign mul_34_17_n_6605 = ~(mul_34_17_n_5324 ^ mul_34_17_n_3093);
 assign mul_34_17_n_6604 = ~(mul_34_17_n_5028 ^ mul_34_17_n_4780);
 assign mul_34_17_n_6602 = ~(mul_34_17_n_5352 ^ mul_34_17_n_2811);
 assign mul_34_17_n_6601 = ~(mul_34_17_n_5284 ^ mul_34_17_n_4451);
 assign mul_34_17_n_6418 = ~(mul_34_17_n_5471 ^ mul_34_17_n_3085);
 assign mul_34_17_n_6417 = (mul_34_17_n_139 ^ mul_34_17_n_4065);
 assign mul_34_17_n_6600 = ~(mul_34_17_n_5472 ^ mul_34_17_n_4748);
 assign mul_34_17_n_6416 = ~(mul_34_17_n_5475 ^ mul_34_17_n_4589);
 assign mul_34_17_n_6599 = ~(mul_34_17_n_5313 ^ mul_34_17_n_4533);
 assign mul_34_17_n_6597 = ~(mul_34_17_n_5280 ^ mul_34_17_n_4677);
 assign mul_34_17_n_6595 = ~(mul_34_17_n_5335 ^ mul_34_17_n_3946);
 assign mul_34_17_n_6594 = ~(mul_34_17_n_5336 ^ mul_34_17_n_4119);
 assign mul_34_17_n_6593 = ~(mul_34_17_n_5343 ^ mul_34_17_n_4765);
 assign mul_34_17_n_6591 = ~(mul_34_17_n_5345 ^ mul_34_17_n_3808);
 assign mul_34_17_n_6590 = ~(mul_34_17_n_5274 ^ mul_34_17_n_4351);
 assign mul_34_17_n_6589 = ~(mul_34_17_n_5273 ^ mul_34_17_n_4344);
 assign mul_34_17_n_6588 = ~(mul_34_17_n_5269 ^ mul_34_17_n_3250);
 assign mul_34_17_n_6586 = ~(mul_34_17_n_5226 ^ mul_34_17_n_4856);
 assign mul_34_17_n_6585 = ~(mul_34_17_n_5268 ^ mul_34_17_n_4580);
 assign mul_34_17_n_6584 = ~(mul_34_17_n_5347 ^ mul_34_17_n_4395);
 assign mul_34_17_n_6581 = ~(mul_34_17_n_5348 ^ mul_34_17_n_4781);
 assign mul_34_17_n_6415 = (mul_34_17_n_5460 ^ mul_34_17_n_4664);
 assign mul_34_17_n_6414 = ~(mul_34_17_n_5459 ^ mul_34_17_n_3824);
 assign mul_34_17_n_6579 = ~(mul_34_17_n_5383 ^ mul_34_17_n_3852);
 assign mul_34_17_n_6577 = ~(mul_34_17_n_5222 ^ mul_34_17_n_4638);
 assign mul_34_17_n_6576 = ~(mul_34_17_n_5218 ^ mul_34_17_n_3809);
 assign mul_34_17_n_6575 = ~(mul_34_17_n_5355 ^ mul_34_17_n_4779);
 assign mul_34_17_n_6574 = ~(mul_34_17_n_5299 ^ mul_34_17_n_3344);
 assign mul_34_17_n_6572 = ~(mul_34_17_n_5259 ^ mul_34_17_n_4702);
 assign mul_34_17_n_6571 = ~(mul_34_17_n_5252 ^ mul_34_17_n_4681);
 assign mul_34_17_n_6570 = ~(mul_34_17_n_5251 ^ mul_34_17_n_4720);
 assign mul_34_17_n_6567 = ~(mul_34_17_n_5356 ^ mul_34_17_n_4792);
 assign mul_34_17_n_6566 = ~(mul_34_17_n_5246 ^ mul_34_17_n_3029);
 assign mul_34_17_n_6565 = ~(mul_34_17_n_5359 ^ mul_34_17_n_4796);
 assign mul_34_17_n_6564 = ~(mul_34_17_n_3962 ^ mul_34_17_n_5244);
 assign mul_34_17_n_6563 = ~(mul_34_17_n_5361 ^ mul_34_17_n_4799);
 assign mul_34_17_n_6561 = ~(mul_34_17_n_5241 ^ mul_34_17_n_4657);
 assign mul_34_17_n_6560 = ~(mul_34_17_n_5248 ^ mul_34_17_n_4279);
 assign mul_34_17_n_6559 = ~(mul_34_17_n_5368 ^ mul_34_17_n_4805);
 assign mul_34_17_n_6557 = ~(mul_34_17_n_5235 ^ mul_34_17_n_4189);
 assign mul_34_17_n_6556 = ~(mul_34_17_n_5234 ^ mul_34_17_n_3183);
 assign mul_34_17_n_6554 = ~(mul_34_17_n_5363 ^ mul_34_17_n_4255);
 assign mul_34_17_n_6413 = ~(mul_34_17_n_5458 ^ mul_34_17_n_2853);
 assign mul_34_17_n_6553 = ~(mul_34_17_n_5279 ^ mul_34_17_n_4089);
 assign mul_34_17_n_6552 = ~(mul_34_17_n_5395 ^ mul_34_17_n_4008);
 assign mul_34_17_n_6550 = ~(mul_34_17_n_5232 ^ mul_34_17_n_4175);
 assign mul_34_17_n_6548 = ~(mul_34_17_n_5229 ^ mul_34_17_n_4172);
 assign mul_34_17_n_6547 = (mul_34_17_n_5486 ^ mul_34_17_n_4717);
 assign mul_34_17_n_6546 = ~(mul_34_17_n_5381 ^ mul_34_17_n_3540);
 assign mul_34_17_n_6545 = ~(mul_34_17_n_5456 ^ mul_34_17_n_4582);
 assign mul_34_17_n_6544 = ~(mul_34_17_n_5455 ^ mul_34_17_n_4018);
 assign mul_34_17_n_6543 = ~(mul_34_17_n_5223 ^ mul_34_17_n_4157);
 assign mul_34_17_n_6542 = ~(mul_34_17_n_5316 ^ mul_34_17_n_4503);
 assign mul_34_17_n_6541 = ~(mul_34_17_n_5219 ^ mul_34_17_n_4768);
 assign mul_34_17_n_6540 = ~(mul_34_17_n_5374 ^ mul_34_17_n_3668);
 assign mul_34_17_n_6539 = ~(mul_34_17_n_5220 ^ mul_34_17_n_4075);
 assign mul_34_17_n_6538 = ~(mul_34_17_n_5051 ^ mul_34_17_n_4608);
 assign mul_34_17_n_6537 = ~(mul_34_17_n_5215 ^ mul_34_17_n_4091);
 assign mul_34_17_n_6536 = ~(mul_34_17_n_5217 ^ mul_34_17_n_4347);
 assign mul_34_17_n_6535 = ~(mul_34_17_n_5375 ^ mul_34_17_n_3666);
 assign mul_34_17_n_6534 = ~(mul_34_17_n_5216 ^ mul_34_17_n_3124);
 assign mul_34_17_n_6533 = ~(mul_34_17_n_5004 ^ mul_34_17_n_3343);
 assign mul_34_17_n_6412 = ~(mul_34_17_n_5488 ^ mul_34_17_n_4812);
 assign mul_34_17_n_6532 = ~(mul_34_17_n_5386 ^ mul_34_17_n_3054);
 assign mul_34_17_n_6411 = ~(mul_34_17_n_5491 ^ mul_34_17_n_3095);
 assign mul_34_17_n_6531 = ~(mul_34_17_n_5376 ^ mul_34_17_n_4818);
 assign mul_34_17_n_6530 = ~(mul_34_17_n_5210 ^ mul_34_17_n_4120);
 assign mul_34_17_n_6529 = ~(mul_34_17_n_5207 ^ mul_34_17_n_4600);
 assign mul_34_17_n_6528 = ~(mul_34_17_n_5206 ^ mul_34_17_n_4653);
 assign mul_34_17_n_6527 = (mul_34_17_n_5467 ^ mul_34_17_n_4714);
 assign mul_34_17_n_6526 = ~(mul_34_17_n_5261 ^ mul_34_17_n_4117);
 assign mul_34_17_n_6525 = ~(mul_34_17_n_5277 ^ mul_34_17_n_4821);
 assign mul_34_17_n_6524 = ~(mul_34_17_n_5228 ^ mul_34_17_n_3814);
 assign mul_34_17_n_6523 = (mul_34_17_n_5461 ^ mul_34_17_n_4676);
 assign mul_34_17_n_6522 = ~(mul_34_17_n_5320 ^ mul_34_17_n_4764);
 assign mul_34_17_n_6520 = ~(mul_34_17_n_5224 ^ mul_34_17_n_4160);
 assign mul_34_17_n_6518 = ~(mul_34_17_n_5369 ^ mul_34_17_n_4685);
 assign mul_34_17_n_6517 = ~(mul_34_17_n_5253 ^ mul_34_17_n_4399);
 assign mul_34_17_n_6516 = ~(mul_34_17_n_5483 ^ mul_34_17_n_4788);
 assign mul_34_17_n_6514 = ~(mul_34_17_n_4988 ^ mul_34_17_n_4552);
 assign mul_34_17_n_6513 = ~(mul_34_17_n_5318 ^ mul_34_17_n_4308);
 assign mul_34_17_n_6511 = ~(mul_34_17_n_5367 ^ mul_34_17_n_4807);
 assign mul_34_17_n_6510 = ~(mul_34_17_n_5302 ^ mul_34_17_n_4159);
 assign mul_34_17_n_6509 = (mul_34_17_n_5169 ^ mul_34_17_n_4619);
 assign mul_34_17_n_6508 = ((mul_34_17_n_4848 & mul_34_17_n_5443) | ((mul_34_17_n_4848 & mul_34_17_n_3561)
    | (mul_34_17_n_3561 & mul_34_17_n_5443)));
 assign mul_34_17_n_6507 = ~(mul_34_17_n_5267 ^ mul_34_17_n_3293);
 assign mul_34_17_n_6506 = ~(mul_34_17_n_5477 ^ mul_34_17_n_4775);
 assign mul_34_17_n_6505 = ~(mul_34_17_n_4998 ^ mul_34_17_n_4123);
 assign mul_34_17_n_6504 = ~(mul_34_17_n_5239 ^ mul_34_17_n_4858);
 assign mul_34_17_n_6503 = ~(mul_34_17_n_5360 ^ mul_34_17_n_4060);
 assign mul_34_17_n_6502 = ~(mul_34_17_n_5480 ^ mul_34_17_n_4789);
 assign mul_34_17_n_6501 = ~(mul_34_17_n_5281 ^ mul_34_17_n_4587);
 assign mul_34_17_n_6500 = ~(mul_34_17_n_5209 ^ mul_34_17_n_3781);
 assign mul_34_17_n_6499 = (mul_34_17_n_5493 ^ mul_34_17_n_4187);
 assign mul_34_17_n_6498 = ~(mul_34_17_n_5365 ^ mul_34_17_n_4802);
 assign mul_34_17_n_6497 = ((mul_34_17_n_3234 & mul_34_17_n_5440) | ((mul_34_17_n_3234 & mul_34_17_n_3235)
    | (mul_34_17_n_3235 & mul_34_17_n_5440)));
 assign mul_34_17_n_6495 = (mul_34_17_n_5453 ^ mul_34_17_n_4620);
 assign mul_34_17_n_6492 = ~(mul_34_17_n_5245 ^ mul_34_17_n_4225);
 assign mul_34_17_n_6489 = ~(mul_34_17_n_5258 ^ mul_34_17_n_4488);
 assign mul_34_17_n_6488 = (mul_34_17_n_5468 ^ mul_34_17_n_4246);
 assign mul_34_17_n_6487 = ~(mul_34_17_n_5272 ^ mul_34_17_n_4397);
 assign mul_34_17_n_6484 = ~(mul_34_17_n_5275 ^ mul_34_17_n_4055);
 assign mul_34_17_n_6483 = ~(mul_34_17_n_5278 ^ mul_34_17_n_4806);
 assign mul_34_17_n_6482 = ~(mul_34_17_n_5462 ^ mul_34_17_n_3591);
 assign mul_34_17_n_6481 = ~(mul_34_17_n_5282 ^ mul_34_17_n_4816);
 assign mul_34_17_n_6480 = ~(mul_34_17_n_4966 ^ mul_34_17_n_4520);
 assign mul_34_17_n_6479 = ~(mul_34_17_n_5283 ^ mul_34_17_n_4705);
 assign mul_34_17_n_6478 = ~(mul_34_17_n_5344 ^ mul_34_17_n_4486);
 assign mul_34_17_n_6477 = ~(mul_34_17_n_5303 ^ mul_34_17_n_4899);
 assign mul_34_17_n_6474 = ~(mul_34_17_n_5305 ^ mul_34_17_n_4740);
 assign mul_34_17_n_6472 = ~(mul_34_17_n_5308 ^ mul_34_17_n_4744);
 assign mul_34_17_n_6471 = ~(mul_34_17_n_5300 ^ mul_34_17_n_4862);
 assign mul_34_17_n_6469 = ~(mul_34_17_n_5319 ^ mul_34_17_n_4762);
 assign mul_34_17_n_6467 = ~(mul_34_17_n_5321 ^ mul_34_17_n_3427);
 assign mul_34_17_n_6466 = ~(mul_34_17_n_5290 ^ mul_34_17_n_3914);
 assign mul_34_17_n_6465 = (mul_34_17_n_5474 ^ mul_34_17_n_4753);
 assign mul_34_17_n_6464 = ~(mul_34_17_n_5479 ^ mul_34_17_n_3691);
 assign mul_34_17_n_6462 = ~(mul_34_17_n_5353 ^ mul_34_17_n_4782);
 assign mul_34_17_n_6461 = ~(mul_34_17_n_5481 ^ mul_34_17_n_2837);
 assign mul_34_17_n_6460 = ~(mul_34_17_n_5484 ^ mul_34_17_n_4791);
 assign mul_34_17_n_6459 = ~(mul_34_17_n_5358 ^ mul_34_17_n_4002);
 assign mul_34_17_n_6458 = ~(mul_34_17_n_5364 ^ mul_34_17_n_4151);
 assign mul_34_17_n_6457 = (mul_34_17_n_5487 ^ mul_34_17_n_4401);
 assign mul_34_17_n_6454 = ((mul_34_17_n_3140 & mul_34_17_n_5450) | ((mul_34_17_n_3140 & mul_34_17_n_3366)
    | (mul_34_17_n_3366 & mul_34_17_n_5450)));
 assign mul_34_17_n_6452 = ~(mul_34_17_n_5208 ^ mul_34_17_n_4607);
 assign mul_34_17_n_6409 = ~mul_34_17_n_6;
 assign mul_34_17_n_6407 = ~mul_34_17_n_6408;
 assign mul_34_17_n_6397 = ~mul_34_17_n_6396;
 assign mul_34_17_n_6393 = ~mul_34_17_n_6392;
 assign mul_34_17_n_6377 = ~mul_34_17_n_6376;
 assign mul_34_17_n_6363 = ~mul_34_17_n_6362;
 assign mul_34_17_n_6353 = ~mul_34_17_n_6352;
 assign mul_34_17_n_6351 = ~mul_34_17_n_6350;
 assign mul_34_17_n_6328 = ~mul_34_17_n_6327;
 assign mul_34_17_n_6308 = ~mul_34_17_n_6309;
 assign mul_34_17_n_6304 = ~mul_34_17_n_6305;
 assign mul_34_17_n_6301 = ~mul_34_17_n_6300;
 assign mul_34_17_n_6299 = ~mul_34_17_n_27;
 assign mul_34_17_n_6269 = ~mul_34_17_n_6268;
 assign mul_34_17_n_6252 = ~mul_34_17_n_6251;
 assign mul_34_17_n_6233 = ~mul_34_17_n_6232;
 assign mul_34_17_n_6231 = ~mul_34_17_n_6230;
 assign mul_34_17_n_6217 = ~mul_34_17_n_6216;
 assign mul_34_17_n_6199 = ~mul_34_17_n_6200;
 assign mul_34_17_n_6193 = ~mul_34_17_n_6194;
 assign mul_34_17_n_6185 = ~mul_34_17_n_6186;
 assign mul_34_17_n_6184 = ~mul_34_17_n_6183;
 assign mul_34_17_n_6177 = ~mul_34_17_n_6178;
 assign mul_34_17_n_6173 = ~mul_34_17_n_6172;
 assign mul_34_17_n_6170 = ~mul_34_17_n_6171;
 assign mul_34_17_n_6152 = ~(mul_34_17_n_5134 ^ mul_34_17_n_3057);
 assign mul_34_17_n_6408 = ~(mul_34_17_n_3967 ^ (mul_34_17_n_4049 ^ (mul_34_17_n_4389 ^ mul_34_17_n_3026)));
 assign mul_34_17_n_6406 = ~(mul_34_17_n_5139 ^ mul_34_17_n_3983);
 assign mul_34_17_n_6147 = (mul_34_17_n_5442 ^ mul_34_17_n_3491);
 assign mul_34_17_n_6405 = ~(mul_34_17_n_5139 ^ mul_34_17_n_3984);
 assign mul_34_17_n_6404 = ~((mul_34_17_n_4390 & mul_34_17_n_3026) | (mul_34_17_n_5203 & mul_34_17_n_77));
 assign mul_34_17_n_6403 = ~(mul_34_17_n_5025 ^ mul_34_17_n_2846);
 assign mul_34_17_n_6402 = ~(mul_34_17_n_5172 ^ mul_34_17_n_3874);
 assign mul_34_17_n_6146 = (mul_34_17_n_5447 ^ mul_34_17_n_4040);
 assign mul_34_17_n_6401 = (mul_34_17_n_5127 ^ mul_34_17_n_3071);
 assign mul_34_17_n_6145 = (mul_34_17_n_4870 ^ mul_34_17_n_5454);
 assign mul_34_17_n_6400 = ~(mul_34_17_n_4927 ^ mul_34_17_n_3704);
 assign mul_34_17_n_6144 = ~(mul_34_17_n_5151 ^ mul_34_17_n_3715);
 assign mul_34_17_n_6399 = ~(mul_34_17_n_4929 ^ mul_34_17_n_3707);
 assign mul_34_17_n_6143 = ~(mul_34_17_n_5150 ^ mul_34_17_n_3208);
 assign mul_34_17_n_6398 = ~(mul_34_17_n_5391 ^ mul_34_17_n_4570);
 assign mul_34_17_n_6396 = ~(mul_34_17_n_5007 ^ mul_34_17_n_4032);
 assign mul_34_17_n_6395 = ~(mul_34_17_n_5121 ^ mul_34_17_n_3065);
 assign mul_34_17_n_6142 = ~(mul_34_17_n_5198 ^ mul_34_17_n_3838);
 assign mul_34_17_n_6394 = ~(mul_34_17_n_5086 ^ mul_34_17_n_3304);
 assign mul_34_17_n_6392 = ~(mul_34_17_n_5080 ^ mul_34_17_n_3738);
 assign mul_34_17_n_6391 = ~(mul_34_17_n_5011 ^ mul_34_17_n_4873);
 assign mul_34_17_n_6141 = (mul_34_17_n_5156 ^ mul_34_17_n_3800);
 assign mul_34_17_n_6390 = ~(mul_34_17_n_5138 ^ mul_34_17_n_3056);
 assign mul_34_17_n_6389 = ~(mul_34_17_n_4960 ^ mul_34_17_n_3807);
 assign mul_34_17_n_6388 = ~(mul_34_17_n_5078 ^ mul_34_17_n_3719);
 assign mul_34_17_n_6387 = ~(mul_34_17_n_4965 ^ mul_34_17_n_3032);
 assign mul_34_17_n_6385 = ~(mul_34_17_n_5075 ^ mul_34_17_n_4066);
 assign mul_34_17_n_6384 = ~(mul_34_17_n_5497 ^ mul_34_17_n_4574);
 assign mul_34_17_n_6382 = ~(mul_34_17_n_4974 ^ mul_34_17_n_3855);
 assign mul_34_17_n_6140 = (mul_34_17_n_5165 ^ mul_34_17_n_3823);
 assign mul_34_17_n_6381 = ~(mul_34_17_n_4980 ^ mul_34_17_n_4640);
 assign mul_34_17_n_6380 = ~(mul_34_17_n_4979 ^ mul_34_17_n_3580);
 assign mul_34_17_n_6379 = ~(mul_34_17_n_4983 ^ mul_34_17_n_4650);
 assign mul_34_17_n_6376 = ~(mul_34_17_n_5044 ^ mul_34_17_n_3689);
 assign mul_34_17_n_6375 = ~(mul_34_17_n_5024 ^ mul_34_17_n_3749);
 assign mul_34_17_n_6374 = ~(mul_34_17_n_4989 ^ mul_34_17_n_4319);
 assign mul_34_17_n_6373 = ~(mul_34_17_n_4992 ^ mul_34_17_n_3760);
 assign mul_34_17_n_6371 = ~(mul_34_17_n_4995 ^ mul_34_17_n_4662);
 assign mul_34_17_n_6370 = ~(mul_34_17_n_4908 ^ mul_34_17_n_3266);
 assign mul_34_17_n_6369 = ~(mul_34_17_n_5066 ^ mul_34_17_n_4794);
 assign mul_34_17_n_6368 = ~(mul_34_17_n_5013 ^ mul_34_17_n_3566);
 assign mul_34_17_n_6139 = ~(mul_34_17_n_5144 ^ mul_34_17_n_2813);
 assign mul_34_17_n_6367 = ~(mul_34_17_n_4917 ^ mul_34_17_n_3168);
 assign mul_34_17_n_6366 = ~(mul_34_17_n_4951 ^ mul_34_17_n_3605);
 assign mul_34_17_n_6365 = ~(mul_34_17_n_5062 ^ mul_34_17_n_3866);
 assign mul_34_17_n_6364 = ~(mul_34_17_n_5331 ^ mul_34_17_n_3034);
 assign mul_34_17_n_6362 = ~(mul_34_17_n_5131 ^ mul_34_17_n_4846);
 assign mul_34_17_n_6361 = ~(mul_34_17_n_4918 ^ mul_34_17_n_3690);
 assign mul_34_17_n_6360 = ~(mul_34_17_n_5037 ^ mul_34_17_n_3786);
 assign mul_34_17_n_6358 = ~(mul_34_17_n_5029 ^ mul_34_17_n_3733);
 assign mul_34_17_n_6357 = ~(mul_34_17_n_5081 ^ mul_34_17_n_3895);
 assign mul_34_17_n_6356 = ~(mul_34_17_n_5130 ^ mul_34_17_n_3976);
 assign mul_34_17_n_6355 = ~(mul_34_17_n_5129 ^ mul_34_17_n_3069);
 assign mul_34_17_n_6354 = ~(mul_34_17_n_5128 ^ mul_34_17_n_3074);
 assign mul_34_17_n_6352 = ~(mul_34_17_n_5047 ^ mul_34_17_n_3903);
 assign mul_34_17_n_6350 = ~(mul_34_17_n_5049 ^ mul_34_17_n_3839);
 assign mul_34_17_n_6138 = (mul_34_17_n_5201 ^ mul_34_17_n_3848);
 assign mul_34_17_n_6349 = ~(mul_34_17_n_5050 ^ mul_34_17_n_3741);
 assign mul_34_17_n_6348 = (mul_34_17_n_5176 ^ mul_34_17_n_4572);
 assign mul_34_17_n_6347 = (mul_34_17_n_5185 ^ mul_34_17_n_3890);
 assign mul_34_17_n_6346 = (mul_34_17_n_5183 ^ mul_34_17_n_4695);
 assign mul_34_17_n_6345 = ~(mul_34_17_n_5182 ^ mul_34_17_n_3900);
 assign mul_34_17_n_6344 = ~(mul_34_17_n_5186 ^ mul_34_17_n_3892);
 assign mul_34_17_n_6343 = ~(mul_34_17_n_5200 ^ mul_34_17_n_4604);
 assign mul_34_17_n_6342 = ~(mul_34_17_n_4948 ^ mul_34_17_n_4847);
 assign mul_34_17_n_6137 = ~(mul_34_17_n_5498 ^ mul_34_17_n_3028);
 assign mul_34_17_n_6341 = ~(mul_34_17_n_5098 ^ mul_34_17_n_3891);
 assign mul_34_17_n_6340 = ~(mul_34_17_n_5043 ^ mul_34_17_n_3734);
 assign mul_34_17_n_6338 = ~(mul_34_17_n_5093 ^ mul_34_17_n_4692);
 assign mul_34_17_n_6336 = ~(mul_34_17_n_5038 ^ mul_34_17_n_3926);
 assign mul_34_17_n_6136 = ~(mul_34_17_n_5187 ^ mul_34_17_n_3879);
 assign mul_34_17_n_6335 = ~(mul_34_17_n_5054 ^ mul_34_17_n_3355);
 assign mul_34_17_n_6334 = ((mul_34_17_n_4355 & mul_34_17_n_5448) | ((mul_34_17_n_4355 & mul_34_17_n_4358)
    | (mul_34_17_n_4358 & mul_34_17_n_5448)));
 assign mul_34_17_n_6333 = ~(mul_34_17_n_5055 ^ mul_34_17_n_3360);
 assign mul_34_17_n_6332 = ~(mul_34_17_n_5298 ^ mul_34_17_n_3869);
 assign mul_34_17_n_6331 = ~(mul_34_17_n_5020 ^ mul_34_17_n_3022);
 assign mul_34_17_n_6330 = (mul_34_17_n_5170 ^ mul_34_17_n_3100);
 assign mul_34_17_n_6329 = (mul_34_17_n_5175 ^ mul_34_17_n_3883);
 assign mul_34_17_n_6327 = ~(mul_34_17_n_5034 ^ mul_34_17_n_3878);
 assign mul_34_17_n_6326 = ~(mul_34_17_n_5392 ^ mul_34_17_n_4003);
 assign mul_34_17_n_6325 = ~(mul_34_17_n_5058 ^ mul_34_17_n_3902);
 assign mul_34_17_n_6324 = ~(mul_34_17_n_5032 ^ mul_34_17_n_3882);
 assign mul_34_17_n_6323 = ~(mul_34_17_n_5056 ^ mul_34_17_n_4254);
 assign mul_34_17_n_6322 = ~(mul_34_17_n_5031 ^ mul_34_17_n_3282);
 assign mul_34_17_n_6320 = ~(mul_34_17_n_5030 ^ mul_34_17_n_3913);
 assign mul_34_17_n_6319 = ~(mul_34_17_n_5059 ^ mul_34_17_n_3739);
 assign mul_34_17_n_6318 = ~(mul_34_17_n_5015 ^ mul_34_17_n_4759);
 assign mul_34_17_n_6317 = ~(mul_34_17_n_5061 ^ mul_34_17_n_3053);
 assign mul_34_17_n_6316 = ~(mul_34_17_n_5026 ^ mul_34_17_n_4605);
 assign mul_34_17_n_6135 = ~(mul_34_17_n_5199 ^ mul_34_17_n_3587);
 assign mul_34_17_n_6315 = ~(mul_34_17_n_5101 ^ mul_34_17_n_4729);
 assign mul_34_17_n_6313 = ~(mul_34_17_n_5385 ^ mul_34_17_n_3583);
 assign mul_34_17_n_6312 = ~(mul_34_17_n_5285 ^ mul_34_17_n_4594);
 assign mul_34_17_n_6311 = ~(mul_34_17_n_5064 ^ mul_34_17_n_3916);
 assign mul_34_17_n_6309 = (mul_34_17_n_5445 ^ mul_34_17_n_2834);
 assign mul_34_17_n_6307 = ~(mul_34_17_n_5018 ^ mul_34_17_n_4869);
 assign mul_34_17_n_6306 = ~(mul_34_17_n_5257 ^ mul_34_17_n_3125);
 assign mul_34_17_n_6305 = ~(mul_34_17_n_5017 ^ mul_34_17_n_4874);
 assign mul_34_17_n_6303 = ~(mul_34_17_n_5191 ^ mul_34_17_n_4700);
 assign mul_34_17_n_6302 = (mul_34_17_n_5192 ^ mul_34_17_n_4691);
 assign mul_34_17_n_6300 = ~(mul_34_17_n_5019 ^ mul_34_17_n_3759);
 assign mul_34_17_n_6134 = (mul_34_17_n_5473 ^ mul_34_17_n_4602);
 assign mul_34_17_n_6298 = ~(mul_34_17_n_5134 ^ mul_34_17_n_3057);
 assign mul_34_17_n_6133 = (mul_34_17_n_5167 ^ mul_34_17_n_4339);
 assign mul_34_17_n_6132 = ~(mul_34_17_n_5166 ^ mul_34_17_n_4001);
 assign mul_34_17_n_6297 = ~(mul_34_17_n_5065 ^ mul_34_17_n_4655);
 assign mul_34_17_n_6296 = ~(mul_34_17_n_5388 ^ mul_34_17_n_4565);
 assign mul_34_17_n_6295 = ~(mul_34_17_n_5000 ^ mul_34_17_n_4643);
 assign mul_34_17_n_6294 = ~(mul_34_17_n_4996 ^ mul_34_17_n_4661);
 assign mul_34_17_n_6291 = ~(mul_34_17_n_5070 ^ mul_34_17_n_2852);
 assign mul_34_17_n_6290 = ~(mul_34_17_n_4993 ^ mul_34_17_n_4312);
 assign mul_34_17_n_6289 = ~(mul_34_17_n_4991 ^ mul_34_17_n_3237);
 assign mul_34_17_n_6287 = ~(mul_34_17_n_4990 ^ mul_34_17_n_4330);
 assign mul_34_17_n_6286 = ~(mul_34_17_n_4938 ^ mul_34_17_n_4688);
 assign mul_34_17_n_6285 = ~(mul_34_17_n_4986 ^ mul_34_17_n_3518);
 assign mul_34_17_n_6284 = ~(mul_34_17_n_4985 ^ mul_34_17_n_3796);
 assign mul_34_17_n_6283 = ~(mul_34_17_n_4984 ^ mul_34_17_n_4642);
 assign mul_34_17_n_6282 = ~(mul_34_17_n_5393 ^ mul_34_17_n_4400);
 assign mul_34_17_n_6281 = ~(mul_34_17_n_4982 ^ mul_34_17_n_4636);
 assign mul_34_17_n_6280 = ~(mul_34_17_n_4981 ^ mul_34_17_n_4861);
 assign mul_34_17_n_6278 = ~(mul_34_17_n_5003 ^ mul_34_17_n_4595);
 assign mul_34_17_n_6277 = ~(mul_34_17_n_5072 ^ mul_34_17_n_3030);
 assign mul_34_17_n_6275 = ~(mul_34_17_n_4973 ^ mul_34_17_n_3437);
 assign mul_34_17_n_6273 = ~(mul_34_17_n_4977 ^ mul_34_17_n_3439);
 assign mul_34_17_n_6271 = ~(mul_34_17_n_4976 ^ mul_34_17_n_3871);
 assign mul_34_17_n_6270 = ~(mul_34_17_n_5090 ^ mul_34_17_n_3428);
 assign mul_34_17_n_6268 = ~(mul_34_17_n_5097 ^ mul_34_17_n_3923);
 assign mul_34_17_n_6267 = ~(mul_34_17_n_4971 ^ mul_34_17_n_3464);
 assign mul_34_17_n_6131 = (mul_34_17_n_5180 ^ mul_34_17_n_4590);
 assign mul_34_17_n_6266 = ~(mul_34_17_n_4969 ^ mul_34_17_n_3468);
 assign mul_34_17_n_6265 = (mul_34_17_n_5184 ^ mul_34_17_n_3886);
 assign mul_34_17_n_6262 = (mul_34_17_n_5164 ^ mul_34_17_n_3780);
 assign mul_34_17_n_6261 = (mul_34_17_n_5163 ^ mul_34_17_n_3777);
 assign mul_34_17_n_6260 = ~(mul_34_17_n_4962 ^ mul_34_17_n_4900);
 assign mul_34_17_n_6259 = ~(mul_34_17_n_5076 ^ mul_34_17_n_3854);
 assign mul_34_17_n_6256 = ~(mul_34_17_n_4959 ^ mul_34_17_n_3412);
 assign mul_34_17_n_6255 = ~(mul_34_17_n_4978 ^ mul_34_17_n_3083);
 assign mul_34_17_n_6254 = ~(mul_34_17_n_5077 ^ mul_34_17_n_3671);
 assign mul_34_17_n_6253 = ~(mul_34_17_n_4955 ^ mul_34_17_n_3768);
 assign mul_34_17_n_6251 = ~(mul_34_17_n_4956 ^ mul_34_17_n_3430);
 assign mul_34_17_n_6250 = ~(mul_34_17_n_4957 ^ mul_34_17_n_4474);
 assign mul_34_17_n_6249 = ~(mul_34_17_n_5099 ^ mul_34_17_n_4808);
 assign mul_34_17_n_6130 = ~(mul_34_17_n_5157 ^ mul_34_17_n_3763);
 assign mul_34_17_n_6248 = ~(mul_34_17_n_5195 ^ mul_34_17_n_3850);
 assign mul_34_17_n_6247 = ~(mul_34_17_n_5153 ^ mul_34_17_n_3764);
 assign mul_34_17_n_6246 = ~(mul_34_17_n_4950 ^ mul_34_17_n_4441);
 assign mul_34_17_n_6245 = ~(mul_34_17_n_4949 ^ mul_34_17_n_3742);
 assign mul_34_17_n_6244 = ~(mul_34_17_n_5196 ^ mul_34_17_n_3722);
 assign mul_34_17_n_6243 = ~(mul_34_17_n_4941 ^ mul_34_17_n_3154);
 assign mul_34_17_n_6242 = ~(mul_34_17_n_4946 ^ mul_34_17_n_3436);
 assign mul_34_17_n_6241 = ~(mul_34_17_n_4945 ^ mul_34_17_n_4860);
 assign mul_34_17_n_6240 = ~(mul_34_17_n_4936 ^ mul_34_17_n_3231);
 assign mul_34_17_n_6239 = ~(mul_34_17_n_5035 ^ mul_34_17_n_3922);
 assign mul_34_17_n_6237 = ~(mul_34_17_n_5247 ^ mul_34_17_n_4368);
 assign mul_34_17_n_6236 = ~(mul_34_17_n_5082 ^ mul_34_17_n_5450);
 assign mul_34_17_n_6235 = ~(mul_34_17_n_4935 ^ mul_34_17_n_3720);
 assign mul_34_17_n_6234 = ~(mul_34_17_n_4915 ^ mul_34_17_n_4154);
 assign mul_34_17_n_6129 = (mul_34_17_n_5171 ^ mul_34_17_n_4865);
 assign mul_34_17_n_6232 = ~(mul_34_17_n_4934 ^ mul_34_17_n_3216);
 assign mul_34_17_n_6230 = ~(mul_34_17_n_5357 ^ mul_34_17_n_3834);
 assign mul_34_17_n_6229 = ~(mul_34_17_n_4910 ^ mul_34_17_n_4262);
 assign mul_34_17_n_6228 = ~(mul_34_17_n_4931 ^ mul_34_17_n_3712);
 assign mul_34_17_n_6227 = ~(mul_34_17_n_5022 ^ mul_34_17_n_3735);
 assign mul_34_17_n_6128 = (mul_34_17_n_5155 ^ mul_34_17_n_3910);
 assign mul_34_17_n_6226 = ~(mul_34_17_n_5088 ^ mul_34_17_n_3826);
 assign mul_34_17_n_6127 = (mul_34_17_n_4864 ^ mul_34_17_n_5149);
 assign mul_34_17_n_6126 = (mul_34_17_n_5148 ^ mul_34_17_n_4571);
 assign mul_34_17_n_6225 = ~(mul_34_17_n_4926 ^ mul_34_17_n_3190);
 assign mul_34_17_n_6224 = ~(mul_34_17_n_5089 ^ mul_34_17_n_3055);
 assign mul_34_17_n_6223 = ~(mul_34_17_n_4914 ^ mul_34_17_n_3182);
 assign mul_34_17_n_6222 = ~(mul_34_17_n_5147 ^ mul_34_17_n_3138);
 assign mul_34_17_n_6221 = ~(mul_34_17_n_4921 ^ mul_34_17_n_3703);
 assign mul_34_17_n_6220 = ~(mul_34_17_n_5146 ^ mul_34_17_n_3697);
 assign mul_34_17_n_6219 = ~(mul_34_17_n_4909 ^ mul_34_17_n_4135);
 assign mul_34_17_n_6125 = (mul_34_17_n_5145 ^ mul_34_17_n_3880);
 assign mul_34_17_n_6218 = (mul_34_17_n_5143 ^ mul_34_17_n_4857);
 assign mul_34_17_n_6216 = ~(mul_34_17_n_5094 ^ mul_34_17_n_4161);
 assign mul_34_17_n_6215 = ~(mul_34_17_n_5095 ^ mul_34_17_n_3911);
 assign mul_34_17_n_6214 = ~(mul_34_17_n_4919 ^ mul_34_17_n_4760);
 assign mul_34_17_n_6213 = ~(mul_34_17_n_5188 ^ mul_34_17_n_3731);
 assign mul_34_17_n_6212 = ~(mul_34_17_n_5085 ^ mul_34_17_n_4697);
 assign mul_34_17_n_6211 = ~(mul_34_17_n_5197 ^ mul_34_17_n_3828);
 assign mul_34_17_n_6210 = ~(mul_34_17_n_4944 ^ mul_34_17_n_4852);
 assign mul_34_17_n_6209 = ~(mul_34_17_n_5159 ^ mul_34_17_n_3767);
 assign mul_34_17_n_6208 = ~(mul_34_17_n_5160 ^ mul_34_17_n_3770);
 assign mul_34_17_n_6206 = ~(mul_34_17_n_4958 ^ mul_34_17_n_3769);
 assign mul_34_17_n_6205 = ~(mul_34_17_n_4967 ^ mul_34_17_n_3139);
 assign mul_34_17_n_6204 = ~(mul_34_17_n_4970 ^ mul_34_17_n_3453);
 assign mul_34_17_n_6203 = ~(mul_34_17_n_4975 ^ mul_34_17_n_2826);
 assign mul_34_17_n_6202 = ~(mul_34_17_n_5194 ^ mul_34_17_n_3920);
 assign mul_34_17_n_6201 = ~(mul_34_17_n_5005 ^ mul_34_17_n_4853);
 assign mul_34_17_n_6200 = (mul_34_17_n_5193 ^ mul_34_17_n_4699);
 assign mul_34_17_n_6198 = ~(mul_34_17_n_5057 ^ mul_34_17_n_4678);
 assign mul_34_17_n_6197 = (mul_34_17_n_5179 ^ mul_34_17_n_3846);
 assign mul_34_17_n_6196 = ~(mul_34_17_n_5496 ^ mul_34_17_n_3615);
 assign mul_34_17_n_6195 = (mul_34_17_n_5482 ^ mul_34_17_n_3745);
 assign mul_34_17_n_6194 = ~(mul_34_17_n_5053 ^ mul_34_17_n_4651);
 assign mul_34_17_n_6192 = ~(mul_34_17_n_5046 ^ mul_34_17_n_4599);
 assign mul_34_17_n_6191 = ~(mul_34_17_n_4923 ^ mul_34_17_n_3771);
 assign mul_34_17_n_6190 = (mul_34_17_n_5178 ^ mul_34_17_n_3686);
 assign mul_34_17_n_6189 = ~(mul_34_17_n_4968 ^ mul_34_17_n_3489);
 assign mul_34_17_n_6188 = ~(mul_34_17_n_4999 ^ mul_34_17_n_3693);
 assign mul_34_17_n_6186 = ~(mul_34_17_n_5039 ^ mul_34_17_n_3862);
 assign mul_34_17_n_6183 = ~(mul_34_17_n_4940 ^ mul_34_17_n_3279);
 assign mul_34_17_n_6182 = (mul_34_17_n_5189 ^ mul_34_17_n_3670);
 assign mul_34_17_n_6181 = ~(mul_34_17_n_4961 ^ mul_34_17_n_3765);
 assign mul_34_17_n_6179 = (mul_34_17_n_5190 ^ mul_34_17_n_3552);
 assign mul_34_17_n_6178 = ~(mul_34_17_n_4939 ^ mul_34_17_n_3724);
 assign mul_34_17_n_6176 = ~(mul_34_17_n_4912 ^ mul_34_17_n_3549);
 assign mul_34_17_n_6175 = ~(mul_34_17_n_4911 ^ mul_34_17_n_4863);
 assign mul_34_17_n_6174 = ~(mul_34_17_n_5067 ^ mul_34_17_n_3756);
 assign mul_34_17_n_6172 = ~(mul_34_17_n_4994 ^ mul_34_17_n_4348);
 assign mul_34_17_n_6171 = ~(mul_34_17_n_5084 ^ mul_34_17_n_4693);
 assign mul_34_17_n_6169 = (mul_34_17_n_5181 ^ mul_34_17_n_4690);
 assign mul_34_17_n_6168 = ~(mul_34_17_n_5168 ^ mul_34_17_n_3805);
 assign mul_34_17_n_6167 = ~(mul_34_17_n_5174 ^ mul_34_17_n_3897);
 assign mul_34_17_n_6166 = (mul_34_17_n_5161 ^ mul_34_17_n_3787);
 assign mul_34_17_n_6165 = ~(mul_34_17_n_5162 ^ mul_34_17_n_3418);
 assign mul_34_17_n_6164 = ~(mul_34_17_n_4972 ^ mul_34_17_n_3459);
 assign mul_34_17_n_6163 = ~(mul_34_17_n_5100 ^ mul_34_17_n_4553);
 assign mul_34_17_n_6162 = (mul_34_17_n_5495 ^ mul_34_17_n_3817);
 assign mul_34_17_n_6161 = ~(mul_34_17_n_4954 ^ mul_34_17_n_4854);
 assign mul_34_17_n_6160 = ~(mul_34_17_n_4997 ^ mul_34_17_n_3998);
 assign mul_34_17_n_6159 = ~(mul_34_17_n_5158 ^ mul_34_17_n_3296);
 assign mul_34_17_n_6158 = ~(mul_34_17_n_5063 ^ mul_34_17_n_3723);
 assign mul_34_17_n_6156 = ~(mul_34_17_n_5069 ^ mul_34_17_n_3678);
 assign mul_34_17_n_6155 = (mul_34_17_n_5154 ^ mul_34_17_n_4659);
 assign mul_34_17_n_6154 = ~(mul_34_17_n_4947 ^ mul_34_17_n_3307);
 assign mul_34_17_n_6153 = ~(mul_34_17_n_5052 ^ mul_34_17_n_2830);
 assign mul_34_17_n_6124 = ~mul_34_17_n_5865;
 assign mul_34_17_n_6123 = ~mul_34_17_n_5856;
 assign mul_34_17_n_6122 = ~mul_34_17_n_5846;
 assign mul_34_17_n_6121 = ~mul_34_17_n_5845;
 assign mul_34_17_n_6120 = ~mul_34_17_n_5844;
 assign mul_34_17_n_6119 = ~mul_34_17_n_5839;
 assign mul_34_17_n_6118 = ~mul_34_17_n_5838;
 assign mul_34_17_n_6114 = ~mul_34_17_n_6113;
 assign mul_34_17_n_6110 = ~mul_34_17_n_6109;
 assign mul_34_17_n_6092 = ~mul_34_17_n_6091;
 assign mul_34_17_n_6079 = ~mul_34_17_n_6078;
 assign mul_34_17_n_6077 = ~mul_34_17_n_6076;
 assign mul_34_17_n_6073 = ~mul_34_17_n_6072;
 assign mul_34_17_n_6069 = ~mul_34_17_n_6068;
 assign mul_34_17_n_6061 = ~mul_34_17_n_6060;
 assign mul_34_17_n_6047 = ~mul_34_17_n_6046;
 assign mul_34_17_n_6030 = ~mul_34_17_n_6029;
 assign mul_34_17_n_6013 = ~mul_34_17_n_6012;
 assign mul_34_17_n_6002 = ~mul_34_17_n_6001;
 assign mul_34_17_n_5999 = ~mul_34_17_n_5998;
 assign mul_34_17_n_5997 = ~mul_34_17_n_5996;
 assign mul_34_17_n_5995 = ~mul_34_17_n_5994;
 assign mul_34_17_n_5993 = ~mul_34_17_n_5992;
 assign mul_34_17_n_5991 = ~mul_34_17_n_5990;
 assign mul_34_17_n_5985 = ~mul_34_17_n_5984;
 assign mul_34_17_n_5983 = ~mul_34_17_n_5982;
 assign mul_34_17_n_5980 = ~mul_34_17_n_5979;
 assign mul_34_17_n_5953 = ~mul_34_17_n_5952;
 assign mul_34_17_n_5950 = ~mul_34_17_n_5949;
 assign mul_34_17_n_5937 = ~mul_34_17_n_5938;
 assign mul_34_17_n_5933 = ~mul_34_17_n_5932;
 assign mul_34_17_n_5931 = ~mul_34_17_n_5930;
 assign mul_34_17_n_5927 = ~mul_34_17_n_5928;
 assign mul_34_17_n_5923 = ~mul_34_17_n_5922;
 assign mul_34_17_n_5912 = ~mul_34_17_n_5911;
 assign mul_34_17_n_5906 = ~mul_34_17_n_5905;
 assign mul_34_17_n_5904 = ~mul_34_17_n_5903;
 assign mul_34_17_n_5897 = ~mul_34_17_n_5898;
 assign mul_34_17_n_5895 = ~mul_34_17_n_5894;
 assign mul_34_17_n_5893 = ~mul_34_17_n_5892;
 assign mul_34_17_n_5890 = ~mul_34_17_n_5889;
 assign mul_34_17_n_5885 = ~mul_34_17_n_5886;
 assign mul_34_17_n_5883 = ~mul_34_17_n_5882;
 assign mul_34_17_n_5878 = ~mul_34_17_n_5879;
 assign mul_34_17_n_5876 = ~mul_34_17_n_5875;
 assign mul_34_17_n_5870 = ~mul_34_17_n_5869;
 assign mul_34_17_n_5868 = ~(mul_34_17_n_5126 & mul_34_17_n_3059);
 assign mul_34_17_n_5867 = ~(mul_34_17_n_5437 & mul_34_17_n_3978);
 assign mul_34_17_n_5866 = ~(mul_34_17_n_5437 | mul_34_17_n_3978);
 assign mul_34_17_n_5865 = ~(mul_34_17_n_5131 & mul_34_17_n_4846);
 assign mul_34_17_n_5864 = ~(mul_34_17_n_5173 & mul_34_17_n_4872);
 assign mul_34_17_n_5863 = ~(mul_34_17_n_5434 & mul_34_17_n_3075);
 assign mul_34_17_n_5862 = ~(mul_34_17_n_5434 | mul_34_17_n_3075);
 assign mul_34_17_n_5861 = ~(mul_34_17_n_5426 & mul_34_17_n_3971);
 assign mul_34_17_n_5860 = ~(mul_34_17_n_5426 | mul_34_17_n_3971);
 assign mul_34_17_n_5859 = ~(mul_34_17_n_5435 | mul_34_17_n_3977);
 assign mul_34_17_n_5858 = ~(mul_34_17_n_5421 & mul_34_17_n_3972);
 assign mul_34_17_n_5857 = ~(mul_34_17_n_5421 | mul_34_17_n_3972);
 assign mul_34_17_n_5856 = ~(mul_34_17_n_5131 | mul_34_17_n_4846);
 assign mul_34_17_n_5855 = ~(mul_34_17_n_5110 & mul_34_17_n_3968);
 assign mul_34_17_n_5854 = ~(mul_34_17_n_5110 | mul_34_17_n_3968);
 assign mul_34_17_n_5853 = ~(mul_34_17_n_5419 & mul_34_17_n_3965);
 assign mul_34_17_n_5852 = ~(mul_34_17_n_5419 | mul_34_17_n_3965);
 assign mul_34_17_n_5851 = ~(mul_34_17_n_5124 | mul_34_17_n_4845);
 assign mul_34_17_n_5850 = ~(mul_34_17_n_5124 & mul_34_17_n_4845);
 assign mul_34_17_n_5849 = ~(mul_34_17_n_5128 | mul_34_17_n_3074);
 assign mul_34_17_n_5848 = ~(mul_34_17_n_5128 & mul_34_17_n_3074);
 assign mul_34_17_n_5847 = ~(mul_34_17_n_5138 | mul_34_17_n_3056);
 assign mul_34_17_n_5846 = ~(mul_34_17_n_5438 | mul_34_17_n_3973);
 assign mul_34_17_n_5845 = ~(mul_34_17_n_5438 & mul_34_17_n_3973);
 assign mul_34_17_n_5844 = ~(mul_34_17_n_5173 | mul_34_17_n_4872);
 assign mul_34_17_n_5843 = ~(mul_34_17_n_5129 & mul_34_17_n_3069);
 assign mul_34_17_n_5842 = ~(mul_34_17_n_5129 | mul_34_17_n_3069);
 assign mul_34_17_n_5841 = ~(mul_34_17_n_5130 | mul_34_17_n_3976);
 assign mul_34_17_n_5840 = ~(mul_34_17_n_5172 & mul_34_17_n_3874);
 assign mul_34_17_n_5839 = ~(mul_34_17_n_5172 | mul_34_17_n_3874);
 assign mul_34_17_n_5838 = ~(mul_34_17_n_5203 & mul_34_17_n_77);
 assign mul_34_17_n_6117 = ~(mul_34_17_n_4851 ^ mul_34_17_n_3087);
 assign mul_34_17_n_5836 = ~(mul_34_17_n_5435 & mul_34_17_n_3977);
 assign mul_34_17_n_5835 = ~(mul_34_17_n_5126 | mul_34_17_n_3059);
 assign mul_34_17_n_5834 = ~(mul_34_17_n_5137 & mul_34_17_n_3062);
 assign mul_34_17_n_5833 = (mul_34_17_n_4849 ^ mul_34_17_n_3300);
 assign mul_34_17_n_5832 = ~(mul_34_17_n_5138 & mul_34_17_n_3056);
 assign mul_34_17_n_5831 = ~(mul_34_17_n_5130 & mul_34_17_n_3976);
 assign mul_34_17_n_6116 = (mul_34_17_n_4851 ^ mul_34_17_n_3087);
 assign mul_34_17_n_5830 = ~(mul_34_17_n_5422 & mul_34_17_n_3974);
 assign mul_34_17_n_5829 = ~(mul_34_17_n_5422 | mul_34_17_n_3974);
 assign mul_34_17_n_5828 = ~(mul_34_17_n_5428 & mul_34_17_n_4885);
 assign mul_34_17_n_5827 = ~(mul_34_17_n_5428 | mul_34_17_n_4885);
 assign mul_34_17_n_5826 = ((mul_34_17_n_4461 & mul_34_17_n_3540) | ((mul_34_17_n_4461 & mul_34_17_n_4466)
    | (mul_34_17_n_4466 & mul_34_17_n_3540)));
 assign mul_34_17_n_5825 = ~((mul_34_17_n_4473 | mul_34_17_n_4478) & (mul_34_17_n_4881 | mul_34_17_n_3969));
 assign mul_34_17_n_5824 = ~((mul_34_17_n_4456 | mul_34_17_n_3118) & (mul_34_17_n_4877 | mul_34_17_n_4451));
 assign mul_34_17_n_5823 = ~(mul_34_17_n_5409 & mul_34_17_n_4879);
 assign mul_34_17_n_5822 = ((mul_34_17_n_4343 & mul_34_17_n_3237) | ((mul_34_17_n_4343 & mul_34_17_n_4133)
    | (mul_34_17_n_4133 & mul_34_17_n_3237)));
 assign mul_34_17_n_5821 = ((mul_34_17_n_4333 & mul_34_17_n_4330) | ((mul_34_17_n_4333 & mul_34_17_n_4337)
    | (mul_34_17_n_4337 & mul_34_17_n_4330)));
 assign mul_34_17_n_5820 = ~(mul_34_17_n_5407 & mul_34_17_n_4882);
 assign mul_34_17_n_5819 = ((mul_34_17_n_3940 | mul_34_17_n_3040) & (mul_34_17_n_4878 | mul_34_17_n_4847));
 assign mul_34_17_n_5818 = ((mul_34_17_n_4322 & mul_34_17_n_4319) | ((mul_34_17_n_4322 & mul_34_17_n_4192)
    | (mul_34_17_n_4192 & mul_34_17_n_4319)));
 assign mul_34_17_n_5817 = ((mul_34_17_n_3350 & mul_34_17_n_3208) | ((mul_34_17_n_3350 & mul_34_17_n_3077)
    | (mul_34_17_n_3077 & mul_34_17_n_3208)));
 assign mul_34_17_n_5816 = ~(mul_34_17_n_5436 | mul_34_17_n_3068);
 assign mul_34_17_n_5814 = ~(mul_34_17_n_5436 & mul_34_17_n_3068);
 assign mul_34_17_n_5813 = (mul_34_17_n_4902 ^ mul_34_17_n_3930);
 assign mul_34_17_n_6115 = ~(mul_34_17_n_4868 ^ mul_34_17_n_2944);
 assign mul_34_17_n_5812 = (mul_34_17_n_3512 ^ mul_34_17_n_4897);
 assign mul_34_17_n_5811 = ~(mul_34_17_n_4859 ^ mul_34_17_n_4310);
 assign mul_34_17_n_5810 = (mul_34_17_n_4178 ^ mul_34_17_n_4888);
 assign mul_34_17_n_5809 = ~(mul_34_17_n_4889 ^ mul_34_17_n_3963);
 assign mul_34_17_n_5808 = ((mul_34_17_n_3522 & mul_34_17_n_4591) | ((mul_34_17_n_3522 & mul_34_17_n_4151)
    | (mul_34_17_n_4151 & mul_34_17_n_4591)));
 assign mul_34_17_n_5807 = ((mul_34_17_n_4102 & mul_34_17_n_4800) | ((mul_34_17_n_4102 & mul_34_17_n_4063)
    | (mul_34_17_n_4063 & mul_34_17_n_4800)));
 assign mul_34_17_n_5806 = ((mul_34_17_n_4373 & mul_34_17_n_4795) | ((mul_34_17_n_4373 & mul_34_17_n_4002)
    | (mul_34_17_n_4002 & mul_34_17_n_4795)));
 assign mul_34_17_n_6113 = ((mul_34_17_n_3321 & mul_34_17_n_4773) | ((mul_34_17_n_3321 & mul_34_17_n_4345)
    | (mul_34_17_n_4345 & mul_34_17_n_4773)));
 assign mul_34_17_n_6112 = ((mul_34_17_n_3117 & mul_34_17_n_3673) | ((mul_34_17_n_3117 & mul_34_17_n_3112)
    | (mul_34_17_n_3112 & mul_34_17_n_3673)));
 assign mul_34_17_n_6111 = ((mul_34_17_n_4088 & mul_34_17_n_4652) | ((mul_34_17_n_4088 & mul_34_17_n_4134)
    | (mul_34_17_n_4134 & mul_34_17_n_4652)));
 assign mul_34_17_n_6109 = ((mul_34_17_n_4235 & mul_34_17_n_4818) | ((mul_34_17_n_4235 & mul_34_17_n_4106)
    | (mul_34_17_n_4106 & mul_34_17_n_4818)));
 assign mul_34_17_n_6108 = ((mul_34_17_n_3408 & mul_34_17_n_4860) | ((mul_34_17_n_3408 & mul_34_17_n_3409)
    | (mul_34_17_n_3409 & mul_34_17_n_4860)));
 assign mul_34_17_n_6107 = ((mul_34_17_n_4257 & mul_34_17_n_3808) | ((mul_34_17_n_4257 & mul_34_17_n_4251)
    | (mul_34_17_n_4251 & mul_34_17_n_3808)));
 assign mul_34_17_n_6106 = ((mul_34_17_n_4456 & mul_34_17_n_4451) | ((mul_34_17_n_4456 & mul_34_17_n_3118)
    | (mul_34_17_n_3118 & mul_34_17_n_4451)));
 assign mul_34_17_n_6105 = ((mul_34_17_n_4084 & mul_34_17_n_4657) | ((mul_34_17_n_4084 & mul_34_17_n_4103)
    | (mul_34_17_n_4103 & mul_34_17_n_4657)));
 assign mul_34_17_n_6104 = ((mul_34_17_n_4009 & mul_34_17_n_4733) | ((mul_34_17_n_4009 & mul_34_17_n_2823)
    | (mul_34_17_n_2823 & mul_34_17_n_4733)));
 assign mul_34_17_n_6103 = ((mul_34_17_n_4555 & mul_34_17_n_4739) | ((mul_34_17_n_4555 & mul_34_17_n_2811)
    | (mul_34_17_n_2811 & mul_34_17_n_4739)));
 assign mul_34_17_n_6102 = ((mul_34_17_n_4311 & mul_34_17_n_4859) | ((mul_34_17_n_4311 & mul_34_17_n_3524)
    | (mul_34_17_n_3524 & mul_34_17_n_4859)));
 assign mul_34_17_n_6101 = ((mul_34_17_n_3356 & mul_34_17_n_3741) | ((mul_34_17_n_3356 & mul_34_17_n_3370)
    | (mul_34_17_n_3370 & mul_34_17_n_3741)));
 assign mul_34_17_n_6100 = ((mul_34_17_n_4444 & mul_34_17_n_3977) | ((mul_34_17_n_4444 & mul_34_17_n_4423)
    | (mul_34_17_n_4423 & mul_34_17_n_3977)));
 assign mul_34_17_n_6099 = ((mul_34_17_n_4431 & mul_34_17_n_3834) | ((mul_34_17_n_4431 & mul_34_17_n_4433)
    | (mul_34_17_n_4433 & mul_34_17_n_3834)));
 assign mul_34_17_n_6098 = ((mul_34_17_n_4277 & mul_34_17_n_4866) | ((mul_34_17_n_4277 & mul_34_17_n_4237)
    | (mul_34_17_n_4237 & mul_34_17_n_4866)));
 assign mul_34_17_n_6097 = ((mul_34_17_n_4331 & mul_34_17_n_4586) | ((mul_34_17_n_4331 & mul_34_17_n_3187)
    | (mul_34_17_n_3187 & mul_34_17_n_4586)));
 assign mul_34_17_n_6096 = ((mul_34_17_n_3349 & mul_34_17_n_3207) | ((mul_34_17_n_3349 & mul_34_17_n_3076)
    | (mul_34_17_n_3076 & mul_34_17_n_3207)));
 assign mul_34_17_n_6095 = ((mul_34_17_n_4360 & mul_34_17_n_4676) | ((mul_34_17_n_4360 & mul_34_17_n_4359)
    | (mul_34_17_n_4359 & mul_34_17_n_4676)));
 assign mul_34_17_n_6094 = ((mul_34_17_n_4351 & mul_34_17_n_4672) | ((mul_34_17_n_4351 & mul_34_17_n_4346)
    | (mul_34_17_n_4346 & mul_34_17_n_4672)));
 assign mul_34_17_n_6093 = ((mul_34_17_n_4287 & mul_34_17_n_3914) | ((mul_34_17_n_4287 & mul_34_17_n_3181)
    | (mul_34_17_n_3181 & mul_34_17_n_3914)));
 assign mul_34_17_n_6091 = ((mul_34_17_n_3653 & mul_34_17_n_3887) | ((mul_34_17_n_3653 & mul_34_17_n_4328)
    | (mul_34_17_n_4328 & mul_34_17_n_3887)));
 assign mul_34_17_n_6090 = ((mul_34_17_n_4306 & mul_34_17_n_4855) | ((mul_34_17_n_4306 & mul_34_17_n_4304)
    | (mul_34_17_n_4304 & mul_34_17_n_4855)));
 assign mul_34_17_n_6089 = ((mul_34_17_n_4259 & mul_34_17_n_4653) | ((mul_34_17_n_4259 & mul_34_17_n_4403)
    | (mul_34_17_n_4403 & mul_34_17_n_4653)));
 assign mul_34_17_n_6088 = ((mul_34_17_n_3182 & mul_34_17_n_3173) | ((mul_34_17_n_3182 & mul_34_17_n_3174)
    | (mul_34_17_n_3174 & mul_34_17_n_3173)));
 assign mul_34_17_n_6087 = ((mul_34_17_n_3238 & mul_34_17_n_3825) | ((mul_34_17_n_3238 & mul_34_17_n_3062)
    | (mul_34_17_n_3062 & mul_34_17_n_3825)));
 assign mul_34_17_n_6086 = ((mul_34_17_n_3620 & mul_34_17_n_3804) | ((mul_34_17_n_3620 & mul_34_17_n_3658)
    | (mul_34_17_n_3658 & mul_34_17_n_3804)));
 assign mul_34_17_n_6085 = ((mul_34_17_n_3169 & mul_34_17_n_4667) | ((mul_34_17_n_3169 & mul_34_17_n_3621)
    | (mul_34_17_n_3621 & mul_34_17_n_4667)));
 assign mul_34_17_n_6084 = ((mul_34_17_n_4137 & mul_34_17_n_3921) | ((mul_34_17_n_4137 & mul_34_17_n_3563)
    | (mul_34_17_n_3563 & mul_34_17_n_3921)));
 assign mul_34_17_n_6083 = ((mul_34_17_n_3553 & mul_34_17_n_4640) | ((mul_34_17_n_3553 & mul_34_17_n_4219)
    | (mul_34_17_n_4219 & mul_34_17_n_4640)));
 assign mul_34_17_n_6082 = ((mul_34_17_n_3102 & mul_34_17_n_3923) | ((mul_34_17_n_3102 & mul_34_17_n_3602)
    | (mul_34_17_n_3602 & mul_34_17_n_3923)));
 assign mul_34_17_n_6081 = ((mul_34_17_n_3502 & mul_34_17_n_3807) | ((mul_34_17_n_3502 & mul_34_17_n_3504)
    | (mul_34_17_n_3504 & mul_34_17_n_3807)));
 assign mul_34_17_n_6080 = ((mul_34_17_n_4197 & mul_34_17_n_4861) | ((mul_34_17_n_4197 & mul_34_17_n_4198)
    | (mul_34_17_n_4198 & mul_34_17_n_4861)));
 assign mul_34_17_n_6078 = ((mul_34_17_n_3617 & mul_34_17_n_3888) | ((mul_34_17_n_3617 & mul_34_17_n_3148)
    | (mul_34_17_n_3148 & mul_34_17_n_3888)));
 assign mul_34_17_n_6076 = ((mul_34_17_n_3558 & mul_34_17_n_4694) | ((mul_34_17_n_3558 & mul_34_17_n_4405)
    | (mul_34_17_n_4405 & mul_34_17_n_4694)));
 assign mul_34_17_n_6075 = ((mul_34_17_n_4119 & mul_34_17_n_4755) | ((mul_34_17_n_4119 & mul_34_17_n_4110)
    | (mul_34_17_n_4110 & mul_34_17_n_4755)));
 assign mul_34_17_n_6074 = ~(mul_34_17_n_5500 & mul_34_17_n_4904);
 assign mul_34_17_n_6072 = ((mul_34_17_n_4125 & mul_34_17_n_4612) | ((mul_34_17_n_4125 & mul_34_17_n_3338)
    | (mul_34_17_n_3338 & mul_34_17_n_4612)));
 assign mul_34_17_n_6071 = ((mul_34_17_n_4531 & mul_34_17_n_4732) | ((mul_34_17_n_4531 & mul_34_17_n_4533)
    | (mul_34_17_n_4533 & mul_34_17_n_4732)));
 assign mul_34_17_n_6070 = ((mul_34_17_n_4145 & mul_34_17_n_4618) | ((mul_34_17_n_4145 & mul_34_17_n_4143)
    | (mul_34_17_n_4143 & mul_34_17_n_4618)));
 assign mul_34_17_n_6068 = ((mul_34_17_n_4126 & mul_34_17_n_4613) | ((mul_34_17_n_4126 & mul_34_17_n_4124)
    | (mul_34_17_n_4124 & mul_34_17_n_4613)));
 assign mul_34_17_n_6067 = ((mul_34_17_n_4261 & mul_34_17_n_4870) | ((mul_34_17_n_4261 & mul_34_17_n_4276)
    | (mul_34_17_n_4276 & mul_34_17_n_4870)));
 assign mul_34_17_n_6066 = ((mul_34_17_n_3297 & mul_34_17_n_3728) | ((mul_34_17_n_3297 & mul_34_17_n_4101)
    | (mul_34_17_n_4101 & mul_34_17_n_3728)));
 assign mul_34_17_n_6065 = ((mul_34_17_n_4093 & mul_34_17_n_3980) | ((mul_34_17_n_4093 & mul_34_17_n_4092)
    | (mul_34_17_n_4092 & mul_34_17_n_3980)));
 assign mul_34_17_n_6064 = ((mul_34_17_n_4077 & mul_34_17_n_4626) | ((mul_34_17_n_4077 & mul_34_17_n_4226)
    | (mul_34_17_n_4226 & mul_34_17_n_4626)));
 assign mul_34_17_n_6063 = ((mul_34_17_n_3339 & mul_34_17_n_3768) | ((mul_34_17_n_3339 & mul_34_17_n_3333)
    | (mul_34_17_n_3333 & mul_34_17_n_3768)));
 assign mul_34_17_n_6062 = ((mul_34_17_n_4090 & mul_34_17_n_4752) | ((mul_34_17_n_4090 & mul_34_17_n_4083)
    | (mul_34_17_n_4083 & mul_34_17_n_4752)));
 assign mul_34_17_n_6060 = ((mul_34_17_n_3348 & mul_34_17_n_4808) | ((mul_34_17_n_3348 & mul_34_17_n_3123)
    | (mul_34_17_n_3123 & mul_34_17_n_4808)));
 assign mul_34_17_n_6059 = ((mul_34_17_n_3528 & mul_34_17_n_3863) | ((mul_34_17_n_3528 & mul_34_17_n_4136)
    | (mul_34_17_n_4136 & mul_34_17_n_3863)));
 assign mul_34_17_n_6058 = ((mul_34_17_n_3421 & mul_34_17_n_3069) | ((mul_34_17_n_3421 & mul_34_17_n_3444)
    | (mul_34_17_n_3444 & mul_34_17_n_3069)));
 assign mul_34_17_n_6057 = ((mul_34_17_n_3516 & mul_34_17_n_3811) | ((mul_34_17_n_3516 & mul_34_17_n_3518)
    | (mul_34_17_n_3518 & mul_34_17_n_3811)));
 assign mul_34_17_n_6056 = ((mul_34_17_n_3315 & mul_34_17_n_3845) | ((mul_34_17_n_3315 & mul_34_17_n_3446)
    | (mul_34_17_n_3446 & mul_34_17_n_3845)));
 assign mul_34_17_n_6055 = ((mul_34_17_n_3210 & mul_34_17_n_3873) | ((mul_34_17_n_3210 & mul_34_17_n_3661)
    | (mul_34_17_n_3661 & mul_34_17_n_3873)));
 assign mul_34_17_n_6054 = ((mul_34_17_n_3192 & mul_34_17_n_3717) | ((mul_34_17_n_3192 & mul_34_17_n_3213)
    | (mul_34_17_n_3213 & mul_34_17_n_3717)));
 assign mul_34_17_n_6053 = ((mul_34_17_n_3569 & mul_34_17_n_4794) | ((mul_34_17_n_3569 & mul_34_17_n_3498)
    | (mul_34_17_n_3498 & mul_34_17_n_4794)));
 assign mul_34_17_n_6052 = ((mul_34_17_n_4371 & mul_34_17_n_3790) | ((mul_34_17_n_4371 & mul_34_17_n_2729)
    | (mul_34_17_n_2729 & mul_34_17_n_3790)));
 assign mul_34_17_n_6051 = ((mul_34_17_n_3594 & mul_34_17_n_3826) | ((mul_34_17_n_3594 & mul_34_17_n_3567)
    | (mul_34_17_n_3567 & mul_34_17_n_3826)));
 assign mul_34_17_n_6050 = ((mul_34_17_n_3457 & mul_34_17_n_3839) | ((mul_34_17_n_3457 & mul_34_17_n_3462)
    | (mul_34_17_n_3462 & mul_34_17_n_3839)));
 assign mul_34_17_n_6049 = ((mul_34_17_n_3431 & mul_34_17_n_4603) | ((mul_34_17_n_3431 & mul_34_17_n_3433)
    | (mul_34_17_n_3433 & mul_34_17_n_4603)));
 assign mul_34_17_n_6048 = ((mul_34_17_n_4338 & mul_34_17_n_4709) | ((mul_34_17_n_4338 & mul_34_17_n_2730)
    | (mul_34_17_n_2730 & mul_34_17_n_4709)));
 assign mul_34_17_n_6046 = ((mul_34_17_n_3354 & mul_34_17_n_3730) | ((mul_34_17_n_3354 & mul_34_17_n_3355)
    | (mul_34_17_n_3355 & mul_34_17_n_3730)));
 assign mul_34_17_n_6045 = ((mul_34_17_n_4522 & mul_34_17_n_4726) | ((mul_34_17_n_4522 & mul_34_17_n_4518)
    | (mul_34_17_n_4518 & mul_34_17_n_4726)));
 assign mul_34_17_n_6044 = ((mul_34_17_n_4007 & mul_34_17_n_4570) | ((mul_34_17_n_4007 & mul_34_17_n_4005)
    | (mul_34_17_n_4005 & mul_34_17_n_4570)));
 assign mul_34_17_n_6043 = ((mul_34_17_n_4203 & mul_34_17_n_4647) | ((mul_34_17_n_4203 & mul_34_17_n_4051)
    | (mul_34_17_n_4051 & mul_34_17_n_4647)));
 assign mul_34_17_n_6042 = ((mul_34_17_n_3555 & mul_34_17_n_4853) | ((mul_34_17_n_3555 & mul_34_17_n_3557)
    | (mul_34_17_n_3557 & mul_34_17_n_4853)));
 assign mul_34_17_n_6041 = ((mul_34_17_n_4548 & mul_34_17_n_4756) | ((mul_34_17_n_4548 & mul_34_17_n_4212)
    | (mul_34_17_n_4212 & mul_34_17_n_4756)));
 assign mul_34_17_n_6040 = ((mul_34_17_n_4480 & mul_34_17_n_3978) | ((mul_34_17_n_4480 & mul_34_17_n_4479)
    | (mul_34_17_n_4479 & mul_34_17_n_3978)));
 assign mul_34_17_n_6039 = ((mul_34_17_n_3129 & mul_34_17_n_4845) | ((mul_34_17_n_3129 & mul_34_17_n_4516)
    | (mul_34_17_n_4516 & mul_34_17_n_4845)));
 assign mul_34_17_n_6038 = ((mul_34_17_n_3445 & mul_34_17_n_3065) | ((mul_34_17_n_3445 & mul_34_17_n_4426)
    | (mul_34_17_n_4426 & mul_34_17_n_3065)));
 assign mul_34_17_n_6037 = ((mul_34_17_n_4385 & mul_34_17_n_4682) | ((mul_34_17_n_4385 & mul_34_17_n_4387)
    | (mul_34_17_n_4387 & mul_34_17_n_4682)));
 assign mul_34_17_n_6036 = ((mul_34_17_n_3342 & mul_34_17_n_4862) | ((mul_34_17_n_3342 & mul_34_17_n_3146)
    | (mul_34_17_n_3146 & mul_34_17_n_4862)));
 assign mul_34_17_n_6035 = ((mul_34_17_n_3332 & mul_34_17_n_4671) | ((mul_34_17_n_3332 & mul_34_17_n_4353)
    | (mul_34_17_n_4353 & mul_34_17_n_4671)));
 assign mul_34_17_n_6034 = ((mul_34_17_n_3416 & mul_34_17_n_3905) | ((mul_34_17_n_3416 & mul_34_17_n_3418)
    | (mul_34_17_n_3418 & mul_34_17_n_3905)));
 assign mul_34_17_n_6033 = ((mul_34_17_n_4363 & mul_34_17_n_4707) | ((mul_34_17_n_4363 & mul_34_17_n_4073)
    | (mul_34_17_n_4073 & mul_34_17_n_4707)));
 assign mul_34_17_n_6032 = ((mul_34_17_n_4294 & mul_34_17_n_3852) | ((mul_34_17_n_4294 & mul_34_17_n_3400)
    | (mul_34_17_n_3400 & mul_34_17_n_3852)));
 assign mul_34_17_n_6031 = ((mul_34_17_n_3590 & mul_34_17_n_3858) | ((mul_34_17_n_3590 & mul_34_17_n_3127)
    | (mul_34_17_n_3127 & mul_34_17_n_3858)));
 assign mul_34_17_n_6029 = ((mul_34_17_n_4497 & mul_34_17_n_4788) | ((mul_34_17_n_4497 & mul_34_17_n_4495)
    | (mul_34_17_n_4495 & mul_34_17_n_4788)));
 assign mul_34_17_n_6028 = ((mul_34_17_n_3227 & mul_34_17_n_3716) | ((mul_34_17_n_3227 & mul_34_17_n_3308)
    | (mul_34_17_n_3308 & mul_34_17_n_3716)));
 assign mul_34_17_n_6027 = ((mul_34_17_n_4086 & mul_34_17_n_4790) | ((mul_34_17_n_4086 & mul_34_17_n_4517)
    | (mul_34_17_n_4517 & mul_34_17_n_4790)));
 assign mul_34_17_n_6026 = ((mul_34_17_n_4344 & mul_34_17_n_4670) | ((mul_34_17_n_4344 & mul_34_17_n_4340)
    | (mul_34_17_n_4340 & mul_34_17_n_4670)));
 assign mul_34_17_n_6025 = ~(mul_34_17_n_4901 ^ mul_34_17_n_4831);
 assign mul_34_17_n_6024 = ((mul_34_17_n_3989 & mul_34_17_n_4823) | ((mul_34_17_n_3989 & mul_34_17_n_4541)
    | (mul_34_17_n_4541 & mul_34_17_n_4823)));
 assign mul_34_17_n_6023 = ((mul_34_17_n_4320 & mul_34_17_n_4673) | ((mul_34_17_n_4320 & mul_34_17_n_4323)
    | (mul_34_17_n_4323 & mul_34_17_n_4673)));
 assign mul_34_17_n_6022 = ((mul_34_17_n_4057 & mul_34_17_n_4580) | ((mul_34_17_n_4057 & mul_34_17_n_4325)
    | (mul_34_17_n_4325 & mul_34_17_n_4580)));
 assign mul_34_17_n_6021 = ((mul_34_17_n_4116 & mul_34_17_n_4814) | ((mul_34_17_n_4116 & mul_34_17_n_4076)
    | (mul_34_17_n_4076 & mul_34_17_n_4814)));
 assign mul_34_17_n_6020 = ((mul_34_17_n_3428 & mul_34_17_n_3664) | ((mul_34_17_n_3428 & mul_34_17_n_3086)
    | (mul_34_17_n_3086 & mul_34_17_n_3664)));
 assign mul_34_17_n_6019 = ((mul_34_17_n_4834 & mul_34_17_n_3036) | ((mul_34_17_n_4834 & mul_34_17_n_4833)
    | (mul_34_17_n_4833 & mul_34_17_n_3036)));
 assign mul_34_17_n_6018 = ((mul_34_17_n_4245 & mul_34_17_n_4584) | ((mul_34_17_n_4245 & mul_34_17_n_2842)
    | (mul_34_17_n_2842 & mul_34_17_n_4584)));
 assign mul_34_17_n_6017 = ((mul_34_17_n_3155 & mul_34_17_n_3721) | ((mul_34_17_n_3155 & mul_34_17_n_3655)
    | (mul_34_17_n_3655 & mul_34_17_n_3721)));
 assign mul_34_17_n_6016 = ((mul_34_17_n_4394 & mul_34_17_n_3761) | ((mul_34_17_n_4394 & mul_34_17_n_4395)
    | (mul_34_17_n_4395 & mul_34_17_n_3761)));
 assign mul_34_17_n_6015 = ((mul_34_17_n_4443 & mul_34_17_n_4810) | ((mul_34_17_n_4443 & mul_34_17_n_4401)
    | (mul_34_17_n_4401 & mul_34_17_n_4810)));
 assign mul_34_17_n_6014 = ((mul_34_17_n_3319 & mul_34_17_n_3910) | ((mul_34_17_n_3319 & mul_34_17_n_3255)
    | (mul_34_17_n_3255 & mul_34_17_n_3910)));
 assign mul_34_17_n_6012 = ((mul_34_17_n_4324 & mul_34_17_n_4768) | ((mul_34_17_n_4324 & mul_34_17_n_3257)
    | (mul_34_17_n_3257 & mul_34_17_n_4768)));
 assign mul_34_17_n_6011 = ((mul_34_17_n_4234 & mul_34_17_n_4589) | ((mul_34_17_n_4234 & mul_34_17_n_3600)
    | (mul_34_17_n_3600 & mul_34_17_n_4589)));
 assign mul_34_17_n_6010 = ((mul_34_17_n_4334 & mul_34_17_n_4348) | ((mul_34_17_n_4334 & mul_34_17_n_4244)
    | (mul_34_17_n_4244 & mul_34_17_n_4348)));
 assign mul_34_17_n_6009 = ((mul_34_17_n_3550 & mul_34_17_n_3738) | ((mul_34_17_n_3550 & mul_34_17_n_3585)
    | (mul_34_17_n_3585 & mul_34_17_n_3738)));
 assign mul_34_17_n_6008 = ((mul_34_17_n_4301 & mul_34_17_n_4771) | ((mul_34_17_n_4301 & mul_34_17_n_4308)
    | (mul_34_17_n_4308 & mul_34_17_n_4771)));
 assign mul_34_17_n_6007 = ((mul_34_17_n_4208 & mul_34_17_n_4636) | ((mul_34_17_n_4208 & mul_34_17_n_4210)
    | (mul_34_17_n_4210 & mul_34_17_n_4636)));
 assign mul_34_17_n_6006 = ((mul_34_17_n_4473 & mul_34_17_n_3969) | ((mul_34_17_n_4473 & mul_34_17_n_4478)
    | (mul_34_17_n_4478 & mul_34_17_n_3969)));
 assign mul_34_17_n_6005 = ((mul_34_17_n_4243 & mul_34_17_n_4767) | ((mul_34_17_n_4243 & mul_34_17_n_4042)
    | (mul_34_17_n_4042 & mul_34_17_n_4767)));
 assign mul_34_17_n_6004 = ((mul_34_17_n_3098 & mul_34_17_n_3667) | ((mul_34_17_n_3098 & mul_34_17_n_3096)
    | (mul_34_17_n_3096 & mul_34_17_n_3667)));
 assign mul_34_17_n_6003 = ((mul_34_17_n_3579 & mul_34_17_n_4867) | ((mul_34_17_n_3579 & mul_34_17_n_4422)
    | (mul_34_17_n_4422 & mul_34_17_n_4867)));
 assign mul_34_17_n_6001 = ((mul_34_17_n_4411 & mul_34_17_n_4698) | ((mul_34_17_n_4411 & mul_34_17_n_2840)
    | (mul_34_17_n_2840 & mul_34_17_n_4698)));
 assign mul_34_17_n_6000 = ((mul_34_17_n_4460 & mul_34_17_n_3539) | ((mul_34_17_n_4460 & mul_34_17_n_4465)
    | (mul_34_17_n_4465 & mul_34_17_n_3539)));
 assign mul_34_17_n_5998 = ((mul_34_17_n_3451 & mul_34_17_n_4758) | ((mul_34_17_n_3451 & mul_34_17_n_4195)
    | (mul_34_17_n_4195 & mul_34_17_n_4758)));
 assign mul_34_17_n_5996 = ((mul_34_17_n_4104 & mul_34_17_n_4751) | ((mul_34_17_n_4104 & mul_34_17_n_4148)
    | (mul_34_17_n_4148 & mul_34_17_n_4751)));
 assign mul_34_17_n_5994 = ((mul_34_17_n_4039 & mul_34_17_n_4746) | ((mul_34_17_n_4039 & mul_34_17_n_4058)
    | (mul_34_17_n_4058 & mul_34_17_n_4746)));
 assign mul_34_17_n_5992 = ((mul_34_17_n_3126 & mul_34_17_n_3675) | ((mul_34_17_n_3126 & mul_34_17_n_3122)
    | (mul_34_17_n_3122 & mul_34_17_n_3675)));
 assign mul_34_17_n_5990 = ((mul_34_17_n_4503 & mul_34_17_n_4757) | ((mul_34_17_n_4503 & mul_34_17_n_4543)
    | (mul_34_17_n_4543 & mul_34_17_n_4757)));
 assign mul_34_17_n_5989 = ((mul_34_17_n_3268 & mul_34_17_n_4847) | ((mul_34_17_n_3268 & mul_34_17_n_4464)
    | (mul_34_17_n_4464 & mul_34_17_n_4847)));
 assign mul_34_17_n_5988 = ((mul_34_17_n_3623 & mul_34_17_n_3867) | ((mul_34_17_n_3623 & mul_34_17_n_4066)
    | (mul_34_17_n_4066 & mul_34_17_n_3867)));
 assign mul_34_17_n_5987 = ((mul_34_17_n_3938 & mul_34_17_n_3035) | ((mul_34_17_n_3938 & mul_34_17_n_3944)
    | (mul_34_17_n_3944 & mul_34_17_n_3035)));
 assign mul_34_17_n_5986 = ((mul_34_17_n_4017 & mul_34_17_n_4624) | ((mul_34_17_n_4017 & mul_34_17_n_4056)
    | (mul_34_17_n_4056 & mul_34_17_n_4624)));
 assign mul_34_17_n_5984 = ((mul_34_17_n_3252 & mul_34_17_n_4600) | ((mul_34_17_n_3252 & mul_34_17_n_3253)
    | (mul_34_17_n_3253 & mul_34_17_n_4600)));
 assign mul_34_17_n_5982 = ((mul_34_17_n_4052 & mul_34_17_n_4797) | ((mul_34_17_n_4052 & mul_34_17_n_4060)
    | (mul_34_17_n_4060 & mul_34_17_n_4797)));
 assign mul_34_17_n_5981 = ((mul_34_17_n_4321 & mul_34_17_n_4318) | ((mul_34_17_n_4321 & mul_34_17_n_4191)
    | (mul_34_17_n_4191 & mul_34_17_n_4318)));
 assign mul_34_17_n_5979 = ((mul_34_17_n_3507 & mul_34_17_n_3812) | ((mul_34_17_n_3507 & mul_34_17_n_3344)
    | (mul_34_17_n_3344 & mul_34_17_n_3812)));
 assign mul_34_17_n_5978 = ((mul_34_17_n_4253 & mul_34_17_n_4684) | ((mul_34_17_n_4253 & mul_34_17_n_3275)
    | (mul_34_17_n_3275 & mul_34_17_n_4684)));
 assign mul_34_17_n_5977 = ((mul_34_17_n_4128 & mul_34_17_n_4750) | ((mul_34_17_n_4128 & mul_34_17_n_4154)
    | (mul_34_17_n_4154 & mul_34_17_n_4750)));
 assign mul_34_17_n_5976 = ((mul_34_17_n_3189 & mul_34_17_n_3692) | ((mul_34_17_n_3189 & mul_34_17_n_3223)
    | (mul_34_17_n_3223 & mul_34_17_n_3692)));
 assign mul_34_17_n_5975 = ((mul_34_17_n_4375 & mul_34_17_n_4778) | ((mul_34_17_n_4375 & mul_34_17_n_4041)
    | (mul_34_17_n_4041 & mul_34_17_n_4778)));
 assign mul_34_17_n_5974 = ((mul_34_17_n_3547 & mul_34_17_n_4597) | ((mul_34_17_n_3547 & mul_34_17_n_4091)
    | (mul_34_17_n_4091 & mul_34_17_n_4597)));
 assign mul_34_17_n_5973 = ((mul_34_17_n_4001 & mul_34_17_n_4598) | ((mul_34_17_n_4001 & mul_34_17_n_2851)
    | (mul_34_17_n_2851 & mul_34_17_n_4598)));
 assign mul_34_17_n_5972 = ((mul_34_17_n_4475 & mul_34_17_n_4713) | ((mul_34_17_n_4475 & mul_34_17_n_4469)
    | (mul_34_17_n_4469 & mul_34_17_n_4713)));
 assign mul_34_17_n_5971 = ((mul_34_17_n_4190 & mul_34_17_n_4761) | ((mul_34_17_n_4190 & mul_34_17_n_3194)
    | (mul_34_17_n_3194 & mul_34_17_n_4761)));
 assign mul_34_17_n_5970 = ((mul_34_17_n_4217 & mul_34_17_n_4721) | ((mul_34_17_n_4217 & mul_34_17_n_4274)
    | (mul_34_17_n_4274 & mul_34_17_n_4721)));
 assign mul_34_17_n_5969 = ((mul_34_17_n_4534 & mul_34_17_n_4735) | ((mul_34_17_n_4534 & mul_34_17_n_4532)
    | (mul_34_17_n_4532 & mul_34_17_n_4735)));
 assign mul_34_17_n_5968 = ((mul_34_17_n_4014 & mul_34_17_n_4569) | ((mul_34_17_n_4014 & mul_34_17_n_3028)
    | (mul_34_17_n_3028 & mul_34_17_n_4569)));
 assign mul_34_17_n_5967 = ((mul_34_17_n_4524 & mul_34_17_n_3073) | ((mul_34_17_n_4524 & mul_34_17_n_4550)
    | (mul_34_17_n_4550 & mul_34_17_n_3073)));
 assign mul_34_17_n_5966 = ((mul_34_17_n_4016 & mul_34_17_n_4873) | ((mul_34_17_n_4016 & mul_34_17_n_4045)
    | (mul_34_17_n_4045 & mul_34_17_n_4873)));
 assign mul_34_17_n_5965 = ((mul_34_17_n_4314 & mul_34_17_n_4312) | ((mul_34_17_n_4314 & mul_34_17_n_4021)
    | (mul_34_17_n_4021 & mul_34_17_n_4312)));
 assign mul_34_17_n_5964 = ((mul_34_17_n_4273 & mul_34_17_n_4805) | ((mul_34_17_n_4273 & mul_34_17_n_4549)
    | (mul_34_17_n_4549 & mul_34_17_n_4805)));
 assign mul_34_17_n_5963 = ((mul_34_17_n_4162 & mul_34_17_n_4689) | ((mul_34_17_n_4162 & mul_34_17_n_4050)
    | (mul_34_17_n_4050 & mul_34_17_n_4689)));
 assign mul_34_17_n_5962 = ((mul_34_17_n_3470 & mul_34_17_n_3074) | ((mul_34_17_n_3470 & mul_34_17_n_3340)
    | (mul_34_17_n_3340 & mul_34_17_n_3074)));
 assign mul_34_17_n_5961 = ((mul_34_17_n_3412 & mul_34_17_n_3778) | ((mul_34_17_n_3412 & mul_34_17_n_3413)
    | (mul_34_17_n_3413 & mul_34_17_n_3778)));
 assign mul_34_17_n_5960 = ((mul_34_17_n_4551 & mul_34_17_n_4711) | ((mul_34_17_n_4551 & mul_34_17_n_4032)
    | (mul_34_17_n_4032 & mul_34_17_n_4711)));
 assign mul_34_17_n_5959 = ((mul_34_17_n_3972 & mul_34_17_n_4745) | ((mul_34_17_n_3972 & mul_34_17_n_4046)
    | (mul_34_17_n_4046 & mul_34_17_n_4745)));
 assign mul_34_17_n_5958 = ((mul_34_17_n_3285 & mul_34_17_n_3854) | ((mul_34_17_n_3285 & mul_34_17_n_3288)
    | (mul_34_17_n_3288 & mul_34_17_n_3854)));
 assign mul_34_17_n_5957 = ((mul_34_17_n_3248 & mul_34_17_n_3734) | ((mul_34_17_n_3248 & mul_34_17_n_3262)
    | (mul_34_17_n_3262 & mul_34_17_n_3734)));
 assign mul_34_17_n_5956 = ((mul_34_17_n_4028 & mul_34_17_n_4744) | ((mul_34_17_n_4028 & mul_34_17_n_4033)
    | (mul_34_17_n_4033 & mul_34_17_n_4744)));
 assign mul_34_17_n_5955 = ((mul_34_17_n_3966 & mul_34_17_n_3736) | ((mul_34_17_n_3966 & mul_34_17_n_2742)
    | (mul_34_17_n_2742 & mul_34_17_n_3736)));
 assign mul_34_17_n_5954 = ((mul_34_17_n_3175 & mul_34_17_n_3719) | ((mul_34_17_n_3175 & mul_34_17_n_3185)
    | (mul_34_17_n_3185 & mul_34_17_n_3719)));
 assign mul_34_17_n_5952 = ((mul_34_17_n_3120 & mul_34_17_n_3685) | ((mul_34_17_n_3120 & mul_34_17_n_3219)
    | (mul_34_17_n_3219 & mul_34_17_n_3685)));
 assign mul_34_17_n_5951 = ((mul_34_17_n_3659 & mul_34_17_n_3671) | ((mul_34_17_n_3659 & mul_34_17_n_3149)
    | (mul_34_17_n_3149 & mul_34_17_n_3671)));
 assign mul_34_17_n_5949 = ((mul_34_17_n_3642 & mul_34_17_n_3926) | ((mul_34_17_n_3642 & mul_34_17_n_3652)
    | (mul_34_17_n_3652 & mul_34_17_n_3926)));
 assign mul_34_17_n_5948 = ((mul_34_17_n_3538 & mul_34_17_n_3821) | ((mul_34_17_n_3538 & mul_34_17_n_3549)
    | (mul_34_17_n_3549 & mul_34_17_n_3821)));
 assign mul_34_17_n_5947 = ((mul_34_17_n_4213 & mul_34_17_n_4639) | ((mul_34_17_n_4213 & mul_34_17_n_3962)
    | (mul_34_17_n_3962 & mul_34_17_n_4639)));
 assign mul_34_17_n_5946 = ((mul_34_17_n_3593 & mul_34_17_n_4688) | ((mul_34_17_n_3593 & mul_34_17_n_4138)
    | (mul_34_17_n_4138 & mul_34_17_n_4688)));
 assign mul_34_17_n_5945 = ((mul_34_17_n_4332 & mul_34_17_n_4329) | ((mul_34_17_n_4332 & mul_34_17_n_4336)
    | (mul_34_17_n_4336 & mul_34_17_n_4329)));
 assign mul_34_17_n_5944 = ((mul_34_17_n_4317 & mul_34_17_n_4) | ((mul_34_17_n_4317 & mul_34_17_n_4316)
    | (mul_34_17_n_4316 & mul_34_17_n_4)));
 assign mul_34_17_n_5943 = ((mul_34_17_n_3221 & mul_34_17_n_3754) | ((mul_34_17_n_3221 & mul_34_17_n_3611)
    | (mul_34_17_n_3611 & mul_34_17_n_3754)));
 assign mul_34_17_n_5942 = ((mul_34_17_n_3530 & mul_34_17_n_4658) | ((mul_34_17_n_3530 & mul_34_17_n_4108)
    | (mul_34_17_n_4108 & mul_34_17_n_4658)));
 assign mul_34_17_n_5941 = ((mul_34_17_n_3196 & mul_34_17_n_4666) | ((mul_34_17_n_3196 & mul_34_17_n_2809)
    | (mul_34_17_n_2809 & mul_34_17_n_4666)));
 assign mul_34_17_n_5940 = ((mul_34_17_n_3133 & mul_34_17_n_4595) | ((mul_34_17_n_3133 & mul_34_17_n_3577)
    | (mul_34_17_n_3577 & mul_34_17_n_4595)));
 assign mul_34_17_n_5939 = ((mul_34_17_n_3099 & mul_34_17_n_3674) | ((mul_34_17_n_3099 & mul_34_17_n_3480)
    | (mul_34_17_n_3480 & mul_34_17_n_3674)));
 assign mul_34_17_n_5938 = ((mul_34_17_n_3450 & mul_34_17_n_3843) | ((mul_34_17_n_3450 & mul_34_17_n_3473)
    | (mul_34_17_n_3473 & mul_34_17_n_3843)));
 assign mul_34_17_n_5936 = ((mul_34_17_n_3466 & mul_34_17_n_3903) | ((mul_34_17_n_3466 & mul_34_17_n_3278)
    | (mul_34_17_n_3278 & mul_34_17_n_3903)));
 assign mul_34_17_n_5935 = ((mul_34_17_n_3056 & mul_34_17_n_3803) | ((mul_34_17_n_3056 & mul_34_17_n_3495)
    | (mul_34_17_n_3495 & mul_34_17_n_3803)));
 assign mul_34_17_n_5934 = ((mul_34_17_n_3107 & mul_34_17_n_3906) | ((mul_34_17_n_3107 & mul_34_17_n_3053)
    | (mul_34_17_n_3053 & mul_34_17_n_3906)));
 assign mul_34_17_n_5932 = ((mul_34_17_n_4078 & mul_34_17_n_4719) | ((mul_34_17_n_4078 & mul_34_17_n_4499)
    | (mul_34_17_n_4499 & mul_34_17_n_4719)));
 assign mul_34_17_n_5930 = ((mul_34_17_n_4491 & mul_34_17_n_4718) | ((mul_34_17_n_4491 & mul_34_17_n_4493)
    | (mul_34_17_n_4493 & mul_34_17_n_4718)));
 assign mul_34_17_n_5929 = ((mul_34_17_n_4438 & mul_34_17_n_3735) | ((mul_34_17_n_4438 & mul_34_17_n_4440)
    | (mul_34_17_n_4440 & mul_34_17_n_3735)));
 assign mul_34_17_n_5928 = ((mul_34_17_n_3303 & mul_34_17_n_3694) | ((mul_34_17_n_3303 & mul_34_17_n_3088)
    | (mul_34_17_n_3088 & mul_34_17_n_3694)));
 assign mul_34_17_n_5926 = ((mul_34_17_n_3381 & mul_34_17_n_3882) | ((mul_34_17_n_3381 & mul_34_17_n_3560)
    | (mul_34_17_n_3560 & mul_34_17_n_3882)));
 assign mul_34_17_n_5925 = ((mul_34_17_n_3584 & mul_34_17_n_3731) | ((mul_34_17_n_3584 & mul_34_17_n_3481)
    | (mul_34_17_n_3481 & mul_34_17_n_3731)));
 assign mul_34_17_n_5924 = ((mul_34_17_n_3361 & mul_34_17_n_4651) | ((mul_34_17_n_3361 & mul_34_17_n_3363)
    | (mul_34_17_n_3363 & mul_34_17_n_4651)));
 assign mul_34_17_n_5922 = ((mul_34_17_n_3599 & mul_34_17_n_3891) | ((mul_34_17_n_3599 & mul_34_17_n_3134)
    | (mul_34_17_n_3134 & mul_34_17_n_3891)));
 assign mul_34_17_n_5921 = ((mul_34_17_n_3973 & mul_34_17_n_4809) | ((mul_34_17_n_3973 & mul_34_17_n_4230)
    | (mul_34_17_n_4230 & mul_34_17_n_4809)));
 assign mul_34_17_n_5920 = ((mul_34_17_n_3059 & mul_34_17_n_4675) | ((mul_34_17_n_3059 & mul_34_17_n_3247)
    | (mul_34_17_n_3247 & mul_34_17_n_4675)));
 assign mul_34_17_n_5919 = ((mul_34_17_n_4357 & mul_34_17_n_4590) | ((mul_34_17_n_4357 & mul_34_17_n_4361)
    | (mul_34_17_n_4361 & mul_34_17_n_4590)));
 assign mul_34_17_n_5918 = ((mul_34_17_n_4068 & mul_34_17_n_4648) | ((mul_34_17_n_4068 & mul_34_17_n_3596)
    | (mul_34_17_n_3596 & mul_34_17_n_4648)));
 assign mul_34_17_n_5917 = ((mul_34_17_n_3331 & mul_34_17_n_3749) | ((mul_34_17_n_3331 & mul_34_17_n_4435)
    | (mul_34_17_n_4435 & mul_34_17_n_3749)));
 assign mul_34_17_n_5916 = ((mul_34_17_n_3358 & mul_34_17_n_3786) | ((mul_34_17_n_3358 & mul_34_17_n_3197)
    | (mul_34_17_n_3197 & mul_34_17_n_3786)));
 assign mul_34_17_n_5915 = ((mul_34_17_n_3199 & mul_34_17_n_3879) | ((mul_34_17_n_3199 & mul_34_17_n_3369)
    | (mul_34_17_n_3369 & mul_34_17_n_3879)));
 assign mul_34_17_n_5914 = ((mul_34_17_n_3398 & mul_34_17_n_4780) | ((mul_34_17_n_3398 & mul_34_17_n_3167)
    | (mul_34_17_n_3167 & mul_34_17_n_4780)));
 assign mul_34_17_n_5913 = ((mul_34_17_n_4003 & mul_34_17_n_4567) | ((mul_34_17_n_4003 & mul_34_17_n_4112)
    | (mul_34_17_n_4112 & mul_34_17_n_4567)));
 assign mul_34_17_n_5911 = ((mul_34_17_n_4376 & mul_34_17_n_4817) | ((mul_34_17_n_4376 & mul_34_17_n_4228)
    | (mul_34_17_n_4228 & mul_34_17_n_4817)));
 assign mul_34_17_n_5910 = ((mul_34_17_n_4207 & mul_34_17_n_4649) | ((mul_34_17_n_4207 & mul_34_17_n_4335)
    | (mul_34_17_n_4335 & mul_34_17_n_4649)));
 assign mul_34_17_n_5909 = ((mul_34_17_n_3266 & mul_34_17_n_3840) | ((mul_34_17_n_3266 & mul_34_17_n_4448)
    | (mul_34_17_n_4448 & mul_34_17_n_3840)));
 assign mul_34_17_n_5908 = ((mul_34_17_n_3454 & mul_34_17_n_3909) | ((mul_34_17_n_3454 & mul_34_17_n_4153)
    | (mul_34_17_n_4153 & mul_34_17_n_3909)));
 assign mul_34_17_n_5907 = ((mul_34_17_n_3990 & mul_34_17_n_4686) | ((mul_34_17_n_3990 & mul_34_17_n_4537)
    | (mul_34_17_n_4537 & mul_34_17_n_4686)));
 assign mul_34_17_n_5905 = ((mul_34_17_n_3605 & mul_34_17_n_3875) | ((mul_34_17_n_3605 & mul_34_17_n_4027)
    | (mul_34_17_n_4027 & mul_34_17_n_3875)));
 assign mul_34_17_n_5903 = ((mul_34_17_n_4233 & mul_34_17_n_4807) | ((mul_34_17_n_4233 & mul_34_17_n_4204)
    | (mul_34_17_n_4204 & mul_34_17_n_4807)));
 assign mul_34_17_n_5902 = ((mul_34_17_n_3310 & mul_34_17_n_4606) | ((mul_34_17_n_3310 & mul_34_17_n_4262)
    | (mul_34_17_n_4262 & mul_34_17_n_4606)));
 assign mul_34_17_n_5901 = ((mul_34_17_n_3535 & mul_34_17_n_3756) | ((mul_34_17_n_3535 & mul_34_17_n_3545)
    | (mul_34_17_n_3545 & mul_34_17_n_3756)));
 assign mul_34_17_n_5900 = ((mul_34_17_n_3509 & mul_34_17_n_3901) | ((mul_34_17_n_3509 & mul_34_17_n_3447)
    | (mul_34_17_n_3447 & mul_34_17_n_3901)));
 assign mul_34_17_n_5899 = ((mul_34_17_n_4238 & mul_34_17_n_4644) | ((mul_34_17_n_4238 & mul_34_17_n_2836)
    | (mul_34_17_n_2836 & mul_34_17_n_4644)));
 assign mul_34_17_n_5898 = ((mul_34_17_n_4265 & mul_34_17_n_4874) | ((mul_34_17_n_4265 & mul_34_17_n_3627)
    | (mul_34_17_n_3627 & mul_34_17_n_4874)));
 assign mul_34_17_n_5896 = ((mul_34_17_n_4121 & mul_34_17_n_4610) | ((mul_34_17_n_4121 & mul_34_17_n_4118)
    | (mul_34_17_n_4118 & mul_34_17_n_4610)));
 assign mul_34_17_n_5894 = ((mul_34_17_n_4498 & mul_34_17_n_4811) | ((mul_34_17_n_4498 & mul_34_17_n_4445)
    | (mul_34_17_n_4445 & mul_34_17_n_4811)));
 assign mul_34_17_n_5892 = ((mul_34_17_n_4074 & mul_34_17_n_4627) | ((mul_34_17_n_4074 & mul_34_17_n_4174)
    | (mul_34_17_n_4174 & mul_34_17_n_4627)));
 assign mul_34_17_n_5891 = ((mul_34_17_n_4510 & mul_34_17_n_4723) | ((mul_34_17_n_4510 & mul_34_17_n_3974)
    | (mul_34_17_n_3974 & mul_34_17_n_4723)));
 assign mul_34_17_n_5889 = ((mul_34_17_n_3572 & mul_34_17_n_3832) | ((mul_34_17_n_3572 & mul_34_17_n_4272)
    | (mul_34_17_n_4272 & mul_34_17_n_3832)));
 assign mul_34_17_n_5888 = ((mul_34_17_n_3613 & mul_34_17_n_4869) | ((mul_34_17_n_3613 & mul_34_17_n_3604)
    | (mul_34_17_n_3604 & mul_34_17_n_4869)));
 assign mul_34_17_n_5887 = ((mul_34_17_n_4342 & mul_34_17_n_3236) | ((mul_34_17_n_4342 & mul_34_17_n_4132)
    | (mul_34_17_n_4132 & mul_34_17_n_3236)));
 assign mul_34_17_n_5886 = ((mul_34_17_n_3597 & mul_34_17_n_3853) | ((mul_34_17_n_3597 & mul_34_17_n_3587)
    | (mul_34_17_n_3587 & mul_34_17_n_3853)));
 assign mul_34_17_n_5884 = ((mul_34_17_n_4525 & mul_34_17_n_4789) | ((mul_34_17_n_4525 & mul_34_17_n_2738)
    | (mul_34_17_n_2738 & mul_34_17_n_4789)));
 assign mul_34_17_n_5882 = ((mul_34_17_n_4379 & mul_34_17_n_4759) | ((mul_34_17_n_4379 & mul_34_17_n_3420)
    | (mul_34_17_n_3420 & mul_34_17_n_4759)));
 assign mul_34_17_n_5881 = ((mul_34_17_n_3437 & mul_34_17_n_3775) | ((mul_34_17_n_3437 & mul_34_17_n_3423)
    | (mul_34_17_n_3423 & mul_34_17_n_3775)));
 assign mul_34_17_n_5880 = ((mul_34_17_n_4457 & mul_34_17_n_4858) | ((mul_34_17_n_4457 & mul_34_17_n_4487)
    | (mul_34_17_n_4487 & mul_34_17_n_4858)));
 assign mul_34_17_n_5879 = ((mul_34_17_n_4454 & mul_34_17_n_3067) | ((mul_34_17_n_4454 & mul_34_17_n_3631)
    | (mul_34_17_n_3631 & mul_34_17_n_3067)));
 assign mul_34_17_n_5877 = ((mul_34_17_n_4519 & mul_34_17_n_3912) | ((mul_34_17_n_4519 & mul_34_17_n_3212)
    | (mul_34_17_n_3212 & mul_34_17_n_3912)));
 assign mul_34_17_n_5875 = ((mul_34_17_n_3265 & mul_34_17_n_3744) | ((mul_34_17_n_3265 & mul_34_17_n_3220)
    | (mul_34_17_n_3220 & mul_34_17_n_3744)));
 assign mul_34_17_n_5874 = ((mul_34_17_n_4229 & mul_34_17_n_4786) | ((mul_34_17_n_4229 & mul_34_17_n_2837)
    | (mul_34_17_n_2837 & mul_34_17_n_4786)));
 assign mul_34_17_n_5872 = ((mul_34_17_n_3328 & mul_34_17_n_3872) | ((mul_34_17_n_3328 & mul_34_17_n_3119)
    | (mul_34_17_n_3119 & mul_34_17_n_3872)));
 assign mul_34_17_n_5871 = ((mul_34_17_n_3443 & mul_34_17_n_4659) | ((mul_34_17_n_3443 & mul_34_17_n_4165)
    | (mul_34_17_n_4165 & mul_34_17_n_4659)));
 assign mul_34_17_n_5869 = ((mul_34_17_n_3496 & mul_34_17_n_3866) | ((mul_34_17_n_3496 & mul_34_17_n_3273)
    | (mul_34_17_n_3273 & mul_34_17_n_3866)));
 assign mul_34_17_n_5790 = ~mul_34_17_n_5789;
 assign mul_34_17_n_5788 = ~mul_34_17_n_5787;
 assign mul_34_17_n_5777 = ~mul_34_17_n_5776;
 assign mul_34_17_n_5768 = ~mul_34_17_n_5767;
 assign mul_34_17_n_5734 = ~mul_34_17_n_5733;
 assign mul_34_17_n_5718 = ~mul_34_17_n_5719;
 assign mul_34_17_n_5703 = ~mul_34_17_n_5702;
 assign mul_34_17_n_5696 = ~mul_34_17_n_5695;
 assign mul_34_17_n_5679 = ~mul_34_17_n_5678;
 assign mul_34_17_n_5674 = ~mul_34_17_n_5673;
 assign mul_34_17_n_5669 = ~mul_34_17_n_5668;
 assign mul_34_17_n_5666 = ~mul_34_17_n_5665;
 assign mul_34_17_n_5658 = ~mul_34_17_n_5657;
 assign mul_34_17_n_5656 = ~mul_34_17_n_5655;
 assign mul_34_17_n_5642 = ~mul_34_17_n_5641;
 assign mul_34_17_n_5633 = ~mul_34_17_n_5632;
 assign mul_34_17_n_5619 = ~mul_34_17_n_5618;
 assign mul_34_17_n_5615 = ~mul_34_17_n_5614;
 assign mul_34_17_n_5613 = ~mul_34_17_n_5612;
 assign mul_34_17_n_5604 = ~mul_34_17_n_5603;
 assign mul_34_17_n_5591 = ~mul_34_17_n_5590;
 assign mul_34_17_n_5586 = ~mul_34_17_n_5585;
 assign mul_34_17_n_5582 = ~mul_34_17_n_5581;
 assign mul_34_17_n_5574 = ~mul_34_17_n_5573;
 assign mul_34_17_n_5560 = ~mul_34_17_n_5559;
 assign mul_34_17_n_5534 = ~mul_34_17_n_5533;
 assign mul_34_17_n_5532 = ~mul_34_17_n_5531;
 assign mul_34_17_n_5530 = ~mul_34_17_n_5529;
 assign mul_34_17_n_5528 = ~mul_34_17_n_5527;
 assign mul_34_17_n_5520 = ~mul_34_17_n_5519;
 assign mul_34_17_n_5516 = ~mul_34_17_n_5515;
 assign mul_34_17_n_5512 = ~mul_34_17_n_5513;
 assign mul_34_17_n_5510 = ~mul_34_17_n_5511;
 assign mul_34_17_n_5506 = ~mul_34_17_n_5507;
 assign mul_34_17_n_5503 = ~(mul_34_17_n_4849 ^ mul_34_17_n_3300);
 assign mul_34_17_n_5502 = ((mul_34_17_n_4200 & mul_34_17_n_4803) | ((mul_34_17_n_4200 & mul_34_17_n_4490)
    | (mul_34_17_n_4490 & mul_34_17_n_4803)));
 assign mul_34_17_n_5501 = (mul_34_17_n_4442 ^ mul_34_17_n_4891);
 assign mul_34_17_n_5805 = ((mul_34_17_n_3646 & mul_34_17_n_4701) | ((mul_34_17_n_3646 & mul_34_17_n_3392)
    | (mul_34_17_n_3392 & mul_34_17_n_4701)));
 assign mul_34_17_n_5804 = ((mul_34_17_n_4038 & mul_34_17_n_4592) | ((mul_34_17_n_4038 & mul_34_17_n_4188)
    | (mul_34_17_n_4188 & mul_34_17_n_4592)));
 assign mul_34_17_n_5803 = ((mul_34_17_n_3352 & mul_34_17_n_4863) | ((mul_34_17_n_3352 & mul_34_17_n_3153)
    | (mul_34_17_n_3153 & mul_34_17_n_4863)));
 assign mul_34_17_n_5802 = ((mul_34_17_n_3165 & mul_34_17_n_3690) | ((mul_34_17_n_3165 & mul_34_17_n_3163)
    | (mul_34_17_n_3163 & mul_34_17_n_3690)));
 assign mul_34_17_n_5801 = ((mul_34_17_n_4408 & mul_34_17_n_3703) | ((mul_34_17_n_4408 & mul_34_17_n_3204)
    | (mul_34_17_n_3204 & mul_34_17_n_3703)));
 assign mul_34_17_n_5800 = ((mul_34_17_n_3292 & mul_34_17_n_4852) | ((mul_34_17_n_3292 & mul_34_17_n_3290)
    | (mul_34_17_n_3290 & mul_34_17_n_4852)));
 assign mul_34_17_n_5799 = ((mul_34_17_n_3097 & mul_34_17_n_3075) | ((mul_34_17_n_3097 & mul_34_17_n_3101)
    | (mul_34_17_n_3101 & mul_34_17_n_3075)));
 assign mul_34_17_n_5798 = ((mul_34_17_n_4062 & mul_34_17_n_4899) | ((mul_34_17_n_4062 & mul_34_17_n_4247)
    | (mul_34_17_n_4247 & mul_34_17_n_4899)));
 assign mul_34_17_n_5797 = ((mul_34_17_n_4474 & mul_34_17_n_4703) | ((mul_34_17_n_4474 & mul_34_17_n_2725)
    | (mul_34_17_n_2725 & mul_34_17_n_4703)));
 assign mul_34_17_n_5796 = ((mul_34_17_n_3373 & mul_34_17_n_4728) | ((mul_34_17_n_3373 & mul_34_17_n_3490)
    | (mul_34_17_n_3490 & mul_34_17_n_4728)));
 assign mul_34_17_n_5795 = ((mul_34_17_n_3459 & mul_34_17_n_3792) | ((mul_34_17_n_3459 & mul_34_17_n_2732)
    | (mul_34_17_n_2732 & mul_34_17_n_3792)));
 assign mul_34_17_n_5794 = ((mul_34_17_n_3209 & mul_34_17_n_4777) | ((mul_34_17_n_3209 & mul_34_17_n_2724)
    | (mul_34_17_n_2724 & mul_34_17_n_4777)));
 assign mul_34_17_n_5793 = ((mul_34_17_n_4558 & mul_34_17_n_4563) | ((mul_34_17_n_4558 & mul_34_17_n_4468)
    | (mul_34_17_n_4468 & mul_34_17_n_4563)));
 assign mul_34_17_n_5792 = ((mul_34_17_n_3514 & mul_34_17_n_4871) | ((mul_34_17_n_3514 & mul_34_17_n_4000)
    | (mul_34_17_n_4000 & mul_34_17_n_4871)));
 assign mul_34_17_n_5791 = ((mul_34_17_n_4396 & mul_34_17_n_4812) | ((mul_34_17_n_4396 & mul_34_17_n_4539)
    | (mul_34_17_n_4539 & mul_34_17_n_4812)));
 assign mul_34_17_n_5789 = ((mul_34_17_n_4221 & mul_34_17_n_4781) | ((mul_34_17_n_4221 & mul_34_17_n_4413)
    | (mul_34_17_n_4413 & mul_34_17_n_4781)));
 assign mul_34_17_n_5787 = ((mul_34_17_n_4356 & mul_34_17_n_4774) | ((mul_34_17_n_4356 & mul_34_17_n_4354)
    | (mul_34_17_n_4354 & mul_34_17_n_4774)));
 assign mul_34_17_n_5786 = ((mul_34_17_n_4209 & mul_34_17_n_4804) | ((mul_34_17_n_4209 & mul_34_17_n_4170)
    | (mul_34_17_n_4170 & mul_34_17_n_4804)));
 assign mul_34_17_n_5785 = ((mul_34_17_n_3971 & mul_34_17_n_3820) | ((mul_34_17_n_3971 & mul_34_17_n_4271)
    | (mul_34_17_n_4271 & mul_34_17_n_3820)));
 assign mul_34_17_n_5784 = ((mul_34_17_n_3057 & mul_34_17_n_3857) | ((mul_34_17_n_3057 & mul_34_17_n_2820)
    | (mul_34_17_n_2820 & mul_34_17_n_3857)));
 assign mul_34_17_n_5783 = ((mul_34_17_n_4224 & mul_34_17_n_4765) | ((mul_34_17_n_4224 & mul_34_17_n_4214)
    | (mul_34_17_n_4214 & mul_34_17_n_4765)));
 assign mul_34_17_n_5782 = ((mul_34_17_n_4010 & mul_34_17_n_4742) | ((mul_34_17_n_4010 & mul_34_17_n_4414)
    | (mul_34_17_n_4414 & mul_34_17_n_4742)));
 assign mul_34_17_n_5781 = ((mul_34_17_n_3105 & mul_34_17_n_3898) | ((mul_34_17_n_3105 & mul_34_17_n_3598)
    | (mul_34_17_n_3598 & mul_34_17_n_3898)));
 assign mul_34_17_n_5780 = ((mul_34_17_n_4546 & mul_34_17_n_4737) | ((mul_34_17_n_4546 & mul_34_17_n_3305)
    | (mul_34_17_n_3305 & mul_34_17_n_4737)));
 assign mul_34_17_n_5779 = ((mul_34_17_n_3280 & mul_34_17_n_3842) | ((mul_34_17_n_3280 & mul_34_17_n_3125)
    | (mul_34_17_n_3125 & mul_34_17_n_3842)));
 assign mul_34_17_n_5778 = ((mul_34_17_n_3091 & mul_34_17_n_3822) | ((mul_34_17_n_3091 & mul_34_17_n_4281)
    | (mul_34_17_n_4281 & mul_34_17_n_3822)));
 assign mul_34_17_n_5776 = ((mul_34_17_n_4507 & mul_34_17_n_4575) | ((mul_34_17_n_4507 & mul_34_17_n_3465)
    | (mul_34_17_n_3465 & mul_34_17_n_4575)));
 assign mul_34_17_n_5775 = ((mul_34_17_n_4485 & mul_34_17_n_4702) | ((mul_34_17_n_4485 & mul_34_17_n_2847)
    | (mul_34_17_n_2847 & mul_34_17_n_4702)));
 assign mul_34_17_n_5774 = ((mul_34_17_n_4449 & mul_34_17_n_4705) | ((mul_34_17_n_4449 & mul_34_17_n_4472)
    | (mul_34_17_n_4472 & mul_34_17_n_4705)));
 assign mul_34_17_n_5773 = ((mul_34_17_n_3131 & mul_34_17_n_4697) | ((mul_34_17_n_3131 & mul_34_17_n_3081)
    | (mul_34_17_n_3081 & mul_34_17_n_4697)));
 assign mul_34_17_n_5772 = ((mul_34_17_n_4072 & mul_34_17_n_4857) | ((mul_34_17_n_4072 & mul_34_17_n_3136)
    | (mul_34_17_n_3136 & mul_34_17_n_4857)));
 assign mul_34_17_n_5771 = ((mul_34_17_n_3570 & mul_34_17_n_3827) | ((mul_34_17_n_3570 & mul_34_17_n_3580)
    | (mul_34_17_n_3580 & mul_34_17_n_3827)));
 assign mul_34_17_n_5770 = ((mul_34_17_n_4377 & mul_34_17_n_4678) | ((mul_34_17_n_4377 & mul_34_17_n_4388)
    | (mul_34_17_n_4388 & mul_34_17_n_4678)));
 assign mul_34_17_n_5769 = ((mul_34_17_n_4381 & mul_34_17_n_4681) | ((mul_34_17_n_4381 & mul_34_17_n_4384)
    | (mul_34_17_n_4384 & mul_34_17_n_4681)));
 assign mul_34_17_n_5767 = ((mul_34_17_n_4169 & mul_34_17_n_4856) | ((mul_34_17_n_4169 & mul_34_17_n_4180)
    | (mul_34_17_n_4180 & mul_34_17_n_4856)));
 assign mul_34_17_n_5766 = ((mul_34_17_n_4299 & mul_34_17_n_3844) | ((mul_34_17_n_4299 & mul_34_17_n_3401)
    | (mul_34_17_n_3401 & mul_34_17_n_3844)));
 assign mul_34_17_n_5765 = ((mul_34_17_n_4285 & mul_34_17_n_3908) | ((mul_34_17_n_4285 & mul_34_17_n_2852)
    | (mul_34_17_n_2852 & mul_34_17_n_3908)));
 assign mul_34_17_n_5764 = ((mul_34_17_n_3484 & mul_34_17_n_4663) | ((mul_34_17_n_3484 & mul_34_17_n_4298)
    | (mul_34_17_n_4298 & mul_34_17_n_4663)));
 assign mul_34_17_n_5763 = ((mul_34_17_n_4218 & mul_34_17_n_4638) | ((mul_34_17_n_4218 & mul_34_17_n_4147)
    | (mul_34_17_n_4147 & mul_34_17_n_4638)));
 assign mul_34_17_n_5762 = ((mul_34_17_n_3402 & mul_34_17_n_4630) | ((mul_34_17_n_3402 & mul_34_17_n_4184)
    | (mul_34_17_n_4184 & mul_34_17_n_4630)));
 assign mul_34_17_n_5761 = ((mul_34_17_n_4043 & mul_34_17_n_3986) | ((mul_34_17_n_4043 & mul_34_17_n_4122)
    | (mul_34_17_n_4122 & mul_34_17_n_3986)));
 assign mul_34_17_n_5760 = ((mul_34_17_n_3083 & mul_34_17_n_4749) | ((mul_34_17_n_3083 & mul_34_17_n_3104)
    | (mul_34_17_n_3104 & mul_34_17_n_4749)));
 assign mul_34_17_n_5759 = ((mul_34_17_n_4283 & mul_34_17_n_4625) | ((mul_34_17_n_4283 & mul_34_17_n_4160)
    | (mul_34_17_n_4160 & mul_34_17_n_4625)));
 assign mul_34_17_n_5758 = ((mul_34_17_n_3394 & mul_34_17_n_4854) | ((mul_34_17_n_3394 & mul_34_17_n_3396)
    | (mul_34_17_n_3396 & mul_34_17_n_4854)));
 assign mul_34_17_n_5757 = ((mul_34_17_n_4374 & mul_34_17_n_4776) | ((mul_34_17_n_4374 & mul_34_17_n_4347)
    | (mul_34_17_n_4347 & mul_34_17_n_4776)));
 assign mul_34_17_n_5756 = ((mul_34_17_n_3525 & mul_34_17_n_3816) | ((mul_34_17_n_3525 & mul_34_17_n_3546)
    | (mul_34_17_n_3546 & mul_34_17_n_3816)));
 assign mul_34_17_n_5755 = ((mul_34_17_n_3240 & mul_34_17_n_3715) | ((mul_34_17_n_3240 & mul_34_17_n_3242)
    | (mul_34_17_n_3242 & mul_34_17_n_3715)));
 assign mul_34_17_n_5754 = ((mul_34_17_n_4189 & mul_34_17_n_4631) | ((mul_34_17_n_4189 & mul_34_17_n_3645)
    | (mul_34_17_n_3645 & mul_34_17_n_4631)));
 assign mul_34_17_n_5753 = ((mul_34_17_n_4095 & mul_34_17_n_4585) | ((mul_34_17_n_4095 & mul_34_17_n_4236)
    | (mul_34_17_n_4236 & mul_34_17_n_4585)));
 assign mul_34_17_n_5752 = ((mul_34_17_n_3657 & mul_34_17_n_4872) | ((mul_34_17_n_3657 & mul_34_17_n_2827)
    | (mul_34_17_n_2827 & mul_34_17_n_4872)));
 assign mul_34_17_n_5751 = ((mul_34_17_n_4182 & mul_34_17_n_4629) | ((mul_34_17_n_4182 & mul_34_17_n_3405)
    | (mul_34_17_n_3405 & mul_34_17_n_4629)));
 assign mul_34_17_n_5750 = ((mul_34_17_n_4020 & mul_34_17_n_3881) | ((mul_34_17_n_4020 & mul_34_17_n_4008)
    | (mul_34_17_n_4008 & mul_34_17_n_3881)));
 assign mul_34_17_n_5749 = ((mul_34_17_n_4047 & mul_34_17_n_4748) | ((mul_34_17_n_4047 & mul_34_17_n_2712)
    | (mul_34_17_n_2712 & mul_34_17_n_4748)));
 assign mul_34_17_n_5748 = ((mul_34_17_n_4462 & mul_34_17_n_4599) | ((mul_34_17_n_4462 & mul_34_17_n_4149)
    | (mul_34_17_n_4149 & mul_34_17_n_4599)));
 assign mul_34_17_n_5747 = ((mul_34_17_n_4542 & mul_34_17_n_4607) | ((mul_34_17_n_4542 & mul_34_17_n_3493)
    | (mul_34_17_n_3493 & mul_34_17_n_4607)));
 assign mul_34_17_n_5746 = ((mul_34_17_n_4378 & mul_34_17_n_4692) | ((mul_34_17_n_4378 & mul_34_17_n_3224)
    | (mul_34_17_n_3224 & mul_34_17_n_4692)));
 assign mul_34_17_n_5745 = ((mul_34_17_n_3404 & mul_34_17_n_4846) | ((mul_34_17_n_3404 & mul_34_17_n_3663)
    | (mul_34_17_n_3663 & mul_34_17_n_4846)));
 assign mul_34_17_n_5744 = ((mul_34_17_n_4284 & mul_34_17_n_3922) | ((mul_34_17_n_4284 & mul_34_17_n_4105)
    | (mul_34_17_n_4105 & mul_34_17_n_3922)));
 assign mul_34_17_n_5743 = ((mul_34_17_n_3618 & mul_34_17_n_3924) | ((mul_34_17_n_3618 & mul_34_17_n_3106)
    | (mul_34_17_n_3106 & mul_34_17_n_3924)));
 assign mul_34_17_n_5742 = ((mul_34_17_n_4196 & mul_34_17_n_4634) | ((mul_34_17_n_4196 & mul_34_17_n_3306)
    | (mul_34_17_n_3306 & mul_34_17_n_4634)));
 assign mul_34_17_n_5741 = ((mul_34_17_n_4225 & mul_34_17_n_4641) | ((mul_34_17_n_4225 & mul_34_17_n_4222)
    | (mul_34_17_n_4222 & mul_34_17_n_4641)));
 assign mul_34_17_n_5740 = ((mul_34_17_n_4111 & mul_34_17_n_4601) | ((mul_34_17_n_4111 & mul_34_17_n_4115)
    | (mul_34_17_n_4115 & mul_34_17_n_4601)));
 assign mul_34_17_n_5739 = ((mul_34_17_n_4267 & mul_34_17_n_3678) | ((mul_34_17_n_4267 & mul_34_17_n_3272)
    | (mul_34_17_n_3272 & mul_34_17_n_3678)));
 assign mul_34_17_n_5738 = ((mul_34_17_n_4064 & mul_34_17_n_3895) | ((mul_34_17_n_4064 & mul_34_17_n_3375)
    | (mul_34_17_n_3375 & mul_34_17_n_3895)));
 assign mul_34_17_n_5737 = ((mul_34_17_n_3193 & mul_34_17_n_4704) | ((mul_34_17_n_3193 & mul_34_17_n_3171)
    | (mul_34_17_n_3171 & mul_34_17_n_4704)));
 assign mul_34_17_n_5736 = ((mul_34_17_n_4459 & mul_34_17_n_3883) | ((mul_34_17_n_4459 & mul_34_17_n_3270)
    | (mul_34_17_n_3270 & mul_34_17_n_3883)));
 assign mul_34_17_n_5735 = ((mul_34_17_n_3619 & mul_34_17_n_3889) | ((mul_34_17_n_3619 & mul_34_17_n_3327)
    | (mul_34_17_n_3327 & mul_34_17_n_3889)));
 assign mul_34_17_n_5733 = ((mul_34_17_n_4263 & mul_34_17_n_4602) | ((mul_34_17_n_4263 & mul_34_17_n_3993)
    | (mul_34_17_n_3993 & mul_34_17_n_4602)));
 assign mul_34_17_n_5732 = ((mul_34_17_n_3186 & mul_34_17_n_4572) | ((mul_34_17_n_3186 & mul_34_17_n_4022)
    | (mul_34_17_n_4022 & mul_34_17_n_4572)));
 assign mul_34_17_n_5731 = ((mul_34_17_n_3565 & mul_34_17_n_3689) | ((mul_34_17_n_3565 & mul_34_17_n_3121)
    | (mul_34_17_n_3121 & mul_34_17_n_3689)));
 assign mul_34_17_n_5730 = ((mul_34_17_n_3371 & mul_34_17_n_3869) | ((mul_34_17_n_3371 & mul_34_17_n_4536)
    | (mul_34_17_n_4536 & mul_34_17_n_3869)));
 assign mul_34_17_n_5729 = ((mul_34_17_n_3510 & mul_34_17_n_3809) | ((mul_34_17_n_3510 & mul_34_17_n_3511)
    | (mul_34_17_n_3511 & mul_34_17_n_3809)));
 assign mul_34_17_n_5728 = ((mul_34_17_n_3474 & mul_34_17_n_3797) | ((mul_34_17_n_3474 & mul_34_17_n_3139)
    | (mul_34_17_n_3139 & mul_34_17_n_3797)));
 assign mul_34_17_n_5727 = ((mul_34_17_n_3458 & mul_34_17_n_3791) | ((mul_34_17_n_3458 & mul_34_17_n_3460)
    | (mul_34_17_n_3460 & mul_34_17_n_3791)));
 assign mul_34_17_n_5726 = ((mul_34_17_n_3410 & mul_34_17_n_3776) | ((mul_34_17_n_3410 & mul_34_17_n_3414)
    | (mul_34_17_n_3414 & mul_34_17_n_3776)));
 assign mul_34_17_n_5725 = ((mul_34_17_n_3374 & mul_34_17_n_3755) | ((mul_34_17_n_3374 & mul_34_17_n_2825)
    | (mul_34_17_n_2825 & mul_34_17_n_3755)));
 assign mul_34_17_n_5724 = ((mul_34_17_n_3382 & mul_34_17_n_3764) | ((mul_34_17_n_3382 & mul_34_17_n_3386)
    | (mul_34_17_n_3386 & mul_34_17_n_3764)));
 assign mul_34_17_n_5723 = ((mul_34_17_n_3378 & mul_34_17_n_3765) | ((mul_34_17_n_3378 & mul_34_17_n_2843)
    | (mul_34_17_n_2843 & mul_34_17_n_3765)));
 assign mul_34_17_n_5722 = ((mul_34_17_n_3161 & mul_34_17_n_3688) | ((mul_34_17_n_3161 & mul_34_17_n_3168)
    | (mul_34_17_n_3168 & mul_34_17_n_3688)));
 assign mul_34_17_n_5721 = ((mul_34_17_n_3286 & mul_34_17_n_4615) | ((mul_34_17_n_3286 & mul_34_17_n_3293)
    | (mul_34_17_n_3293 & mul_34_17_n_4615)));
 assign mul_34_17_n_5720 = ((mul_34_17_n_3316 & mul_34_17_n_3740) | ((mul_34_17_n_3316 & mul_34_17_n_4441)
    | (mul_34_17_n_4441 & mul_34_17_n_3740)));
 assign mul_34_17_n_5719 = ((mul_34_17_n_3461 & mul_34_17_n_3796) | ((mul_34_17_n_3461 & mul_34_17_n_3456)
    | (mul_34_17_n_3456 & mul_34_17_n_3796)));
 assign mul_34_17_n_5717 = ((mul_34_17_n_3222 & mul_34_17_n_3712) | ((mul_34_17_n_3222 & mul_34_17_n_2835)
    | (mul_34_17_n_2835 & mul_34_17_n_3712)));
 assign mul_34_17_n_5716 = ((mul_34_17_n_3274 & mul_34_17_n_3727) | ((mul_34_17_n_3274 & mul_34_17_n_3279)
    | (mul_34_17_n_3279 & mul_34_17_n_3727)));
 assign mul_34_17_n_5715 = ((mul_34_17_n_3322 & mul_34_17_n_3835) | ((mul_34_17_n_3322 & mul_34_17_n_3079)
    | (mul_34_17_n_3079 & mul_34_17_n_3835)));
 assign mul_34_17_n_5714 = ((mul_34_17_n_3492 & mul_34_17_n_3030) | ((mul_34_17_n_3492 & mul_34_17_n_3505)
    | (mul_34_17_n_3505 & mul_34_17_n_3030)));
 assign mul_34_17_n_5713 = ((mul_34_17_n_3997 & mul_34_17_n_4565) | ((mul_34_17_n_3997 & mul_34_17_n_3995)
    | (mul_34_17_n_3995 & mul_34_17_n_4565)));
 assign mul_34_17_n_5712 = ((mul_34_17_n_4425 & mul_34_17_n_4700) | ((mul_34_17_n_4425 & mul_34_17_n_4428)
    | (mul_34_17_n_4428 & mul_34_17_n_4700)));
 assign mul_34_17_n_5711 = ((mul_34_17_n_4419 & mul_34_17_n_4699) | ((mul_34_17_n_4419 & mul_34_17_n_4421)
    | (mul_34_17_n_4421 & mul_34_17_n_4699)));
 assign mul_34_17_n_5710 = ((mul_34_17_n_4250 & mul_34_17_n_3029) | ((mul_34_17_n_4250 & mul_34_17_n_4241)
    | (mul_34_17_n_4241 & mul_34_17_n_3029)));
 assign mul_34_17_n_5709 = ((mul_34_17_n_4398 & mul_34_17_n_4685) | ((mul_34_17_n_4398 & mul_34_17_n_4070)
    | (mul_34_17_n_4070 & mul_34_17_n_4685)));
 assign mul_34_17_n_5708 = ((mul_34_17_n_3337 & mul_34_17_n_3032) | ((mul_34_17_n_3337 & mul_34_17_n_3229)
    | (mul_34_17_n_3229 & mul_34_17_n_3032)));
 assign mul_34_17_n_5707 = ((mul_34_17_n_3425 & mul_34_17_n_4900) | ((mul_34_17_n_3425 & mul_34_17_n_3581)
    | (mul_34_17_n_3581 & mul_34_17_n_4900)));
 assign mul_34_17_n_5706 = ((mul_34_17_n_3232 & mul_34_17_n_3711) | ((mul_34_17_n_3232 & mul_34_17_n_3250)
    | (mul_34_17_n_3250 & mul_34_17_n_3711)));
 assign mul_34_17_n_5705 = ((mul_34_17_n_3142 & mul_34_17_n_4886) | ((mul_34_17_n_3142 & mul_34_17_n_3144)
    | (mul_34_17_n_3144 & mul_34_17_n_4886)));
 assign mul_34_17_n_5704 = ((mul_34_17_n_3641 & mul_34_17_n_3877) | ((mul_34_17_n_3641 & mul_34_17_n_4161)
    | (mul_34_17_n_4161 & mul_34_17_n_3877)));
 assign mul_34_17_n_5702 = ((mul_34_17_n_3372 & mul_34_17_n_3762) | ((mul_34_17_n_3372 & mul_34_17_n_4167)
    | (mul_34_17_n_4167 & mul_34_17_n_3762)));
 assign mul_34_17_n_5701 = ((mul_34_17_n_3998 & mul_34_17_n_3753) | ((mul_34_17_n_3998 & mul_34_17_n_3987)
    | (mul_34_17_n_3987 & mul_34_17_n_3753)));
 assign mul_34_17_n_5700 = ((mul_34_17_n_4553 & mul_34_17_n_3752) | ((mul_34_17_n_4553 & mul_34_17_n_4526)
    | (mul_34_17_n_4526 & mul_34_17_n_3752)));
 assign mul_34_17_n_5699 = ((mul_34_17_n_4268 & mul_34_17_n_4683) | ((mul_34_17_n_4268 & mul_34_17_n_3334)
    | (mul_34_17_n_3334 & mul_34_17_n_4683)));
 assign mul_34_17_n_5698 = ((mul_34_17_n_4365 & mul_34_17_n_4677) | ((mul_34_17_n_4365 & mul_34_17_n_4364)
    | (mul_34_17_n_4364 & mul_34_17_n_4677)));
 assign mul_34_17_n_5697 = ((mul_34_17_n_4146 & mul_34_17_n_4798) | ((mul_34_17_n_4146 & mul_34_17_n_4256)
    | (mul_34_17_n_4256 & mul_34_17_n_4798)));
 assign mul_34_17_n_5695 = ((mul_34_17_n_4307 & mul_34_17_n_3760) | ((mul_34_17_n_4307 & mul_34_17_n_4309)
    | (mul_34_17_n_4309 & mul_34_17_n_3760)));
 assign mul_34_17_n_5694 = ((mul_34_17_n_3326 & mul_34_17_n_3729) | ((mul_34_17_n_3326 & mul_34_17_n_4523)
    | (mul_34_17_n_4523 & mul_34_17_n_3729)));
 assign mul_34_17_n_5693 = ((mul_34_17_n_4291 & mul_34_17_n_4661) | ((mul_34_17_n_4291 & mul_34_17_n_3640)
    | (mul_34_17_n_3640 & mul_34_17_n_4661)));
 assign mul_34_17_n_5692 = ((mul_34_17_n_3320 & mul_34_17_n_4581) | ((mul_34_17_n_3320 & mul_34_17_n_2717)
    | (mul_34_17_n_2717 & mul_34_17_n_4581)));
 assign mul_34_17_n_5691 = ((mul_34_17_n_4352 & mul_34_17_n_4583) | ((mul_34_17_n_4352 & mul_34_17_n_4055)
    | (mul_34_17_n_4055 & mul_34_17_n_4583)));
 assign mul_34_17_n_5690 = ((mul_34_17_n_3455 & mul_34_17_n_3739) | ((mul_34_17_n_3455 & mul_34_17_n_2721)
    | (mul_34_17_n_2721 & mul_34_17_n_3739)));
 assign mul_34_17_n_5689 = ((mul_34_17_n_4297 & mul_34_17_n_3824) | ((mul_34_17_n_4297 & mul_34_17_n_4296)
    | (mul_34_17_n_4296 & mul_34_17_n_3824)));
 assign mul_34_17_n_5688 = ((mul_34_17_n_3092 & mul_34_17_n_3871) | ((mul_34_17_n_3092 & mul_34_17_n_3170)
    | (mul_34_17_n_3170 & mul_34_17_n_3871)));
 assign mul_34_17_n_5687 = ((mul_34_17_n_4127 & mul_34_17_n_4611) | ((mul_34_17_n_4127 & mul_34_17_n_2853)
    | (mul_34_17_n_2853 & mul_34_17_n_4611)));
 assign mul_34_17_n_5686 = ((mul_34_17_n_3654 & mul_34_17_n_3864) | ((mul_34_17_n_3654 & mul_34_17_n_4386)
    | (mul_34_17_n_4386 & mul_34_17_n_3864)));
 assign mul_34_17_n_5685 = ((mul_34_17_n_4249 & mul_34_17_n_4650) | ((mul_34_17_n_4249 & mul_34_17_n_3508)
    | (mul_34_17_n_3508 & mul_34_17_n_4650)));
 assign mul_34_17_n_5684 = ((mul_34_17_n_3629 & mul_34_17_n_3851) | ((mul_34_17_n_3629 & mul_34_17_n_4382)
    | (mul_34_17_n_4382 & mul_34_17_n_3851)));
 assign mul_34_17_n_5683 = ((mul_34_17_n_4471 & mul_34_17_n_4779) | ((mul_34_17_n_4471 & mul_34_17_n_4415)
    | (mul_34_17_n_4415 & mul_34_17_n_4779)));
 assign mul_34_17_n_5682 = ((mul_34_17_n_4227 & mul_34_17_n_4642) | ((mul_34_17_n_4227 & mul_34_17_n_4085)
    | (mul_34_17_n_4085 & mul_34_17_n_4642)));
 assign mul_34_17_n_5681 = ((mul_34_17_n_3566 & mul_34_17_n_3830) | ((mul_34_17_n_3566 & mul_34_17_n_2736)
    | (mul_34_17_n_2736 & mul_34_17_n_3830)));
 assign mul_34_17_n_5680 = ((mul_34_17_n_3159 & mul_34_17_n_3870) | ((mul_34_17_n_3159 & mul_34_17_n_3116)
    | (mul_34_17_n_3116 & mul_34_17_n_3870)));
 assign mul_34_17_n_5678 = ((mul_34_17_n_4406 & mul_34_17_n_3693) | ((mul_34_17_n_4406 & mul_34_17_n_4477)
    | (mul_34_17_n_4477 & mul_34_17_n_3693)));
 assign mul_34_17_n_5677 = ((mul_34_17_n_4201 & mul_34_17_n_4635) | ((mul_34_17_n_4201 & mul_34_17_n_4081)
    | (mul_34_17_n_4081 & mul_34_17_n_4635)));
 assign mul_34_17_n_5676 = ((mul_34_17_n_3531 & mul_34_17_n_3841) | ((mul_34_17_n_3531 & mul_34_17_n_4194)
    | (mul_34_17_n_4194 & mul_34_17_n_3841)));
 assign mul_34_17_n_5675 = ((mul_34_17_n_3520 & mul_34_17_n_3810) | ((mul_34_17_n_3520 & mul_34_17_n_2735)
    | (mul_34_17_n_2735 & mul_34_17_n_3810)));
 assign mul_34_17_n_5673 = ((mul_34_17_n_4141 & mul_34_17_n_3907) | ((mul_34_17_n_4141 & mul_34_17_n_3551)
    | (mul_34_17_n_3551 & mul_34_17_n_3907)));
 assign mul_34_17_n_5672 = ((mul_34_17_n_4031 & mul_34_17_n_4743) | ((mul_34_17_n_4031 & mul_34_17_n_4019)
    | (mul_34_17_n_4019 & mul_34_17_n_4743)));
 assign mul_34_17_n_5671 = ((mul_34_17_n_3215 & mul_34_17_n_3710) | ((mul_34_17_n_3215 & mul_34_17_n_2816)
    | (mul_34_17_n_2816 & mul_34_17_n_3710)));
 assign mul_34_17_n_5670 = ((mul_34_17_n_4561 & mul_34_17_n_4796) | ((mul_34_17_n_4561 & mul_34_17_n_4545)
    | (mul_34_17_n_4545 & mul_34_17_n_4796)));
 assign mul_34_17_n_5668 = ((mul_34_17_n_4175 & mul_34_17_n_3894) | ((mul_34_17_n_4175 & mul_34_17_n_3526)
    | (mul_34_17_n_3526 & mul_34_17_n_3894)));
 assign mul_34_17_n_5667 = ((mul_34_17_n_3203 & mul_34_17_n_4864) | ((mul_34_17_n_3203 & mul_34_17_n_3201)
    | (mul_34_17_n_3201 & mul_34_17_n_4864)));
 assign mul_34_17_n_5665 = ((mul_34_17_n_4368 & mul_34_17_n_3868) | ((mul_34_17_n_4368 & mul_34_17_n_3564)
    | (mul_34_17_n_3564 & mul_34_17_n_3868)));
 assign mul_34_17_n_5664 = ((mul_34_17_n_4144 & mul_34_17_n_3681) | ((mul_34_17_n_4144 & mul_34_17_n_3124)
    | (mul_34_17_n_3124 & mul_34_17_n_3681)));
 assign mul_34_17_n_5663 = ((mul_34_17_n_4173 & mul_34_17_n_4706) | ((mul_34_17_n_4173 & mul_34_17_n_3218)
    | (mul_34_17_n_3218 & mul_34_17_n_4706)));
 assign mul_34_17_n_5662 = ((mul_34_17_n_3230 & mul_34_17_n_3714) | ((mul_34_17_n_3230 & mul_34_17_n_2723)
    | (mul_34_17_n_2723 & mul_34_17_n_3714)));
 assign mul_34_17_n_5661 = ((mul_34_17_n_3137 & mul_34_17_n_3698) | ((mul_34_17_n_3137 & mul_34_17_n_2727)
    | (mul_34_17_n_2727 & mul_34_17_n_3698)));
 assign mul_34_17_n_5660 = ((mul_34_17_n_4075 & mul_34_17_n_4621) | ((mul_34_17_n_4075 & mul_34_17_n_4150)
    | (mul_34_17_n_4150 & mul_34_17_n_4621)));
 assign mul_34_17_n_5659 = ((mul_34_17_n_4193 & mul_34_17_n_4815) | ((mul_34_17_n_4193 & mul_34_17_n_3606)
    | (mul_34_17_n_3606 & mul_34_17_n_4815)));
 assign mul_34_17_n_5657 = ((mul_34_17_n_4107 & mul_34_17_n_4763) | ((mul_34_17_n_4107 & mul_34_17_n_4065)
    | (mul_34_17_n_4065 & mul_34_17_n_4763)));
 assign mul_34_17_n_5655 = ((mul_34_17_n_4131 & mul_34_17_n_3758) | ((mul_34_17_n_4131 & mul_34_17_n_4186)
    | (mul_34_17_n_4186 & mul_34_17_n_3758)));
 assign mul_34_17_n_5654 = ((mul_34_17_n_4447 & mul_34_17_n_4620) | ((mul_34_17_n_4447 & mul_34_17_n_3245)
    | (mul_34_17_n_3245 & mul_34_17_n_4620)));
 assign mul_34_17_n_5653 = ((mul_34_17_n_3307 & mul_34_17_n_3737) | ((mul_34_17_n_3307 & mul_34_17_n_2819)
    | (mul_34_17_n_2819 & mul_34_17_n_3737)));
 assign mul_34_17_n_5652 = ((mul_34_17_n_4292 & mul_34_17_n_4821) | ((mul_34_17_n_4292 & mul_34_17_n_4059)
    | (mul_34_17_n_4059 & mul_34_17_n_4821)));
 assign mul_34_17_n_5651 = ((mul_34_17_n_4130 & mul_34_17_n_4614) | ((mul_34_17_n_4130 & mul_34_17_n_4129)
    | (mul_34_17_n_4129 & mul_34_17_n_4614)));
 assign mul_34_17_n_5650 = ((mul_34_17_n_4482 & mul_34_17_n_4816) | ((mul_34_17_n_4482 & mul_34_17_n_4140)
    | (mul_34_17_n_4140 & mul_34_17_n_4816)));
 assign mul_34_17_n_5649 = ((mul_34_17_n_4290 & mul_34_17_n_4820) | ((mul_34_17_n_4290 & mul_34_17_n_4024)
    | (mul_34_17_n_4024 & mul_34_17_n_4820)));
 assign mul_34_17_n_5648 = ((mul_34_17_n_4183 & mul_34_17_n_3876) | ((mul_34_17_n_4183 & mul_34_17_n_3183)
    | (mul_34_17_n_3183 & mul_34_17_n_3876)));
 assign mul_34_17_n_5647 = ((mul_34_17_n_4171 & mul_34_17_n_4628) | ((mul_34_17_n_4171 & mul_34_17_n_4172)
    | (mul_34_17_n_4172 & mul_34_17_n_4628)));
 assign mul_34_17_n_5646 = ((mul_34_17_n_4206 & mul_34_17_n_4637) | ((mul_34_17_n_4206 & mul_34_17_n_4205)
    | (mul_34_17_n_4205 & mul_34_17_n_4637)));
 assign mul_34_17_n_5645 = ((mul_34_17_n_4362 & mul_34_17_n_4806) | ((mul_34_17_n_4362 & mul_34_17_n_4392)
    | (mul_34_17_n_4392 & mul_34_17_n_4806)));
 assign mul_34_17_n_5644 = ((mul_34_17_n_4254 & mul_34_17_n_4793) | ((mul_34_17_n_4254 & mul_34_17_n_3082)
    | (mul_34_17_n_3082 & mul_34_17_n_4793)));
 assign mul_34_17_n_5643 = ((mul_34_17_n_3992 & mul_34_17_n_4669) | ((mul_34_17_n_3992 & mul_34_17_n_4216)
    | (mul_34_17_n_4216 & mul_34_17_n_4669)));
 assign mul_34_17_n_5641 = ((mul_34_17_n_3506 & mul_34_17_n_3669) | ((mul_34_17_n_3506 & mul_34_17_n_3103)
    | (mul_34_17_n_3103 & mul_34_17_n_3669)));
 assign mul_34_17_n_5640 = ((mul_34_17_n_4452 & mul_34_17_n_3859) | ((mul_34_17_n_4452 & mul_34_17_n_4450)
    | (mul_34_17_n_4450 & mul_34_17_n_3859)));
 assign mul_34_17_n_5639 = ((mul_34_17_n_3548 & mul_34_17_n_3836) | ((mul_34_17_n_3548 & mul_34_17_n_3529)
    | (mul_34_17_n_3529 & mul_34_17_n_3836)));
 assign mul_34_17_n_5638 = ((mul_34_17_n_3486 & mul_34_17_n_3837) | ((mul_34_17_n_3486 & mul_34_17_n_3426)
    | (mul_34_17_n_3426 & mul_34_17_n_3837)));
 assign mul_34_17_n_5637 = ((mul_34_17_n_4407 & mul_34_17_n_4747) | ((mul_34_17_n_4407 & mul_34_17_n_4393)
    | (mul_34_17_n_4393 & mul_34_17_n_4747)));
 assign mul_34_17_n_5636 = ((mul_34_17_n_3991 & mul_34_17_n_4716) | ((mul_34_17_n_3991 & mul_34_17_n_4556)
    | (mul_34_17_n_4556 & mul_34_17_n_4716)));
 assign mul_34_17_n_5635 = ((mul_34_17_n_4114 & mul_34_17_n_3781) | ((mul_34_17_n_4114 & mul_34_17_n_4113)
    | (mul_34_17_n_4113 & mul_34_17_n_3781)));
 assign mul_34_17_n_5634 = ((mul_34_17_n_3313 & mul_34_17_n_3885) | ((mul_34_17_n_3313 & mul_34_17_n_2830)
    | (mul_34_17_n_2830 & mul_34_17_n_3885)));
 assign mul_34_17_n_5632 = ((mul_34_17_n_3314 & mul_34_17_n_3742) | ((mul_34_17_n_3314 & mul_34_17_n_3309)
    | (mul_34_17_n_3309 & mul_34_17_n_3742)));
 assign mul_34_17_n_5631 = ((mul_34_17_n_3628 & mul_34_17_n_3672) | ((mul_34_17_n_3628 & mul_34_17_n_3583)
    | (mul_34_17_n_3583 & mul_34_17_n_3672)));
 assign mul_34_17_n_5630 = ((mul_34_17_n_3055 & mul_34_17_n_4734) | ((mul_34_17_n_3055 & mul_34_17_n_3609)
    | (mul_34_17_n_3609 & mul_34_17_n_4734)));
 assign mul_34_17_n_5629 = ((mul_34_17_n_3357 & mul_34_17_n_3748) | ((mul_34_17_n_3357 & mul_34_17_n_3367)
    | (mul_34_17_n_3367 & mul_34_17_n_3748)));
 assign mul_34_17_n_5628 = ((mul_34_17_n_3284 & mul_34_17_n_3984) | ((mul_34_17_n_3284 & mul_34_17_n_3283)
    | (mul_34_17_n_3283 & mul_34_17_n_3984)));
 assign mul_34_17_n_5627 = ((mul_34_17_n_3467 & mul_34_17_n_3788) | ((mul_34_17_n_3467 & mul_34_17_n_3499)
    | (mul_34_17_n_3499 & mul_34_17_n_3788)));
 assign mul_34_17_n_5626 = ((mul_34_17_n_3260 & mul_34_17_n_3918) | ((mul_34_17_n_3260 & mul_34_17_n_3296)
    | (mul_34_17_n_3296 & mul_34_17_n_3918)));
 assign mul_34_17_n_5625 = ((mul_34_17_n_3312 & mul_34_17_n_3828) | ((mul_34_17_n_3312 & mul_34_17_n_4240)
    | (mul_34_17_n_4240 & mul_34_17_n_3828)));
 assign mul_34_17_n_5624 = ((mul_34_17_n_4370 & mul_34_17_n_3691) | ((mul_34_17_n_4370 & mul_34_17_n_4367)
    | (mul_34_17_n_4367 & mul_34_17_n_3691)));
 assign mul_34_17_n_5623 = ((mul_34_17_n_4053 & mul_34_17_n_4656) | ((mul_34_17_n_4053 & mul_34_17_n_3638)
    | (mul_34_17_n_3638 & mul_34_17_n_4656)));
 assign mul_34_17_n_5622 = ((mul_34_17_n_3616 & mul_34_17_n_3925) | ((mul_34_17_n_3616 & mul_34_17_n_3633)
    | (mul_34_17_n_3633 & mul_34_17_n_3925)));
 assign mul_34_17_n_5621 = ((mul_34_17_n_4527 & mul_34_17_n_4730) | ((mul_34_17_n_4527 & mul_34_17_n_4429)
    | (mul_34_17_n_4429 & mul_34_17_n_4730)));
 assign mul_34_17_n_5620 = ((mul_34_17_n_4069 & mul_34_17_n_3981) | ((mul_34_17_n_4069 & mul_34_17_n_4079)
    | (mul_34_17_n_4079 & mul_34_17_n_3981)));
 assign mul_34_17_n_5618 = ((mul_34_17_n_4269 & mul_34_17_n_4792) | ((mul_34_17_n_4269 & mul_34_17_n_4535)
    | (mul_34_17_n_4535 & mul_34_17_n_4792)));
 assign mul_34_17_n_5617 = ((mul_34_17_n_4098 & mul_34_17_n_4801) | ((mul_34_17_n_4098 & mul_34_17_n_2818)
    | (mul_34_17_n_2818 & mul_34_17_n_4801)));
 assign mul_34_17_n_5616 = ((mul_34_17_n_4313 & mul_34_17_n_4772) | ((mul_34_17_n_4313 & mul_34_17_n_4341)
    | (mul_34_17_n_4341 & mul_34_17_n_4772)));
 assign mul_34_17_n_5614 = ((mul_34_17_n_3586 & mul_34_17_n_3915) | ((mul_34_17_n_3586 & mul_34_17_n_3573)
    | (mul_34_17_n_3573 & mul_34_17_n_3915)));
 assign mul_34_17_n_5612 = ((mul_34_17_n_3406 & mul_34_17_n_3896) | ((mul_34_17_n_3406 & mul_34_17_n_3650)
    | (mul_34_17_n_3650 & mul_34_17_n_3896)));
 assign mul_34_17_n_5611 = ((mul_34_17_n_4538 & mul_34_17_n_4787) | ((mul_34_17_n_4538 & mul_34_17_n_4315)
    | (mul_34_17_n_4315 & mul_34_17_n_4787)));
 assign mul_34_17_n_5610 = ((mul_34_17_n_3376 & mul_34_17_n_3913) | ((mul_34_17_n_3376 & mul_34_17_n_4467)
    | (mul_34_17_n_4467 & mul_34_17_n_3913)));
 assign mul_34_17_n_5609 = ((mul_34_17_n_3543 & mul_34_17_n_3683) | ((mul_34_17_n_3543 & mul_34_17_n_2813)
    | (mul_34_17_n_2813 & mul_34_17_n_3683)));
 assign mul_34_17_n_5608 = ((mul_34_17_n_3536 & mul_34_17_n_3865) | ((mul_34_17_n_3536 & mul_34_17_n_3362)
    | (mul_34_17_n_3362 & mul_34_17_n_3865)));
 assign mul_34_17_n_5607 = ((mul_34_17_n_4232 & mul_34_17_n_4764) | ((mul_34_17_n_4232 & mul_34_17_n_3589)
    | (mul_34_17_n_3589 & mul_34_17_n_4764)));
 assign mul_34_17_n_5606 = ((mul_34_17_n_3287 & mul_34_17_n_3884) | ((mul_34_17_n_3287 & mul_34_17_n_3614)
    | (mul_34_17_n_3614 & mul_34_17_n_3884)));
 assign mul_34_17_n_5605 = ((mul_34_17_n_3276 & mul_34_17_n_4708) | ((mul_34_17_n_3276 & mul_34_17_n_3282)
    | (mul_34_17_n_3282 & mul_34_17_n_4708)));
 assign mul_34_17_n_5603 = ((mul_34_17_n_4402 & mul_34_17_n_3886) | ((mul_34_17_n_4402 & mul_34_17_n_3302)
    | (mul_34_17_n_3302 & mul_34_17_n_3886)));
 assign mul_34_17_n_5602 = ((mul_34_17_n_3441 & mul_34_17_n_4633) | ((mul_34_17_n_3441 & mul_34_17_n_3353)
    | (mul_34_17_n_3353 & mul_34_17_n_4633)));
 assign mul_34_17_n_5601 = ((mul_34_17_n_4455 & mul_34_17_n_4622) | ((mul_34_17_n_4455 & mul_34_17_n_4470)
    | (mul_34_17_n_4470 & mul_34_17_n_4622)));
 assign mul_34_17_n_5600 = ((mul_34_17_n_3347 & mul_34_17_n_3892) | ((mul_34_17_n_3347 & mul_34_17_n_3346)
    | (mul_34_17_n_3346 & mul_34_17_n_3892)));
 assign mul_34_17_n_5599 = ((mul_34_17_n_4417 & mul_34_17_n_4782) | ((mul_34_17_n_4417 & mul_34_17_n_4416)
    | (mul_34_17_n_4416 & mul_34_17_n_4782)));
 assign mul_34_17_n_5598 = ((mul_34_17_n_4026 & mul_34_17_n_4573) | ((mul_34_17_n_4026 & mul_34_17_n_4025)
    | (mul_34_17_n_4025 & mul_34_17_n_4573)));
 assign mul_34_17_n_5597 = ((mul_34_17_n_4012 & mul_34_17_n_4579) | ((mul_34_17_n_4012 & mul_34_17_n_4302)
    | (mul_34_17_n_4302 & mul_34_17_n_4579)));
 assign mul_34_17_n_5596 = ((mul_34_17_n_3154 & mul_34_17_n_3676) | ((mul_34_17_n_3154 & mul_34_17_n_3176)
    | (mul_34_17_n_3176 & mul_34_17_n_3676)));
 assign mul_34_17_n_5595 = ((mul_34_17_n_3054 & mul_34_17_n_4577) | ((mul_34_17_n_3054 & mul_34_17_n_4035)
    | (mul_34_17_n_4035 & mul_34_17_n_4577)));
 assign mul_34_17_n_5594 = ((mul_34_17_n_3562 & mul_34_17_n_3829) | ((mul_34_17_n_3562 & mul_34_17_n_3323)
    | (mul_34_17_n_3323 & mul_34_17_n_3829)));
 assign mul_34_17_n_5593 = ((mul_34_17_n_4258 & mul_34_17_n_4660) | ((mul_34_17_n_4258 & mul_34_17_n_3147)
    | (mul_34_17_n_3147 & mul_34_17_n_4660)));
 assign mul_34_17_n_5592 = ((mul_34_17_n_3637 & mul_34_17_n_3916) | ((mul_34_17_n_3637 & mul_34_17_n_3647)
    | (mul_34_17_n_3647 & mul_34_17_n_3916)));
 assign mul_34_17_n_5590 = ((mul_34_17_n_3377 & mul_34_17_n_3766) | ((mul_34_17_n_3377 & mul_34_17_n_3379)
    | (mul_34_17_n_3379 & mul_34_17_n_3766)));
 assign mul_34_17_n_5589 = ((mul_34_17_n_4559 & mul_34_17_n_4587) | ((mul_34_17_n_4559 & mul_34_17_n_4547)
    | (mul_34_17_n_4547 & mul_34_17_n_4587)));
 assign mul_34_17_n_5588 = ((mul_34_17_n_3335 & mul_34_17_n_3070) | ((mul_34_17_n_3335 & mul_34_17_n_4061)
    | (mul_34_17_n_4061 & mul_34_17_n_3070)));
 assign mul_34_17_n_5587 = ((mul_34_17_n_3111 & mul_34_17_n_3757) | ((mul_34_17_n_3111 & mul_34_17_n_3094)
    | (mul_34_17_n_3094 & mul_34_17_n_3757)));
 assign mul_34_17_n_5585 = ((mul_34_17_n_3258 & mul_34_17_n_4632) | ((mul_34_17_n_3258 & mul_34_17_n_4120)
    | (mul_34_17_n_4120 & mul_34_17_n_4632)));
 assign mul_34_17_n_5584 = ((mul_34_17_n_3150 & mul_34_17_n_3861) | ((mul_34_17_n_3150 & mul_34_17_n_2849)
    | (mul_34_17_n_2849 & mul_34_17_n_3861)));
 assign mul_34_17_n_5583 = ((mul_34_17_n_3533 & mul_34_17_n_3818) | ((mul_34_17_n_3533 & mul_34_17_n_3537)
    | (mul_34_17_n_3537 & mul_34_17_n_3818)));
 assign mul_34_17_n_5581 = ((mul_34_17_n_3517 & mul_34_17_n_3814) | ((mul_34_17_n_3517 & mul_34_17_n_3521)
    | (mul_34_17_n_3521 & mul_34_17_n_3814)));
 assign mul_34_17_n_5580 = ((mul_34_17_n_4544 & mul_34_17_n_4729) | ((mul_34_17_n_4544 & mul_34_17_n_4554)
    | (mul_34_17_n_4554 & mul_34_17_n_4729)));
 assign mul_34_17_n_5579 = ((mul_34_17_n_3294 & mul_34_17_n_4645) | ((mul_34_17_n_3294 & mul_34_17_n_4279)
    | (mul_34_17_n_4279 & mul_34_17_n_4645)));
 assign mul_34_17_n_5578 = ((mul_34_17_n_3299 & mul_34_17_n_3849) | ((mul_34_17_n_3299 & mul_34_17_n_3295)
    | (mul_34_17_n_3295 & mul_34_17_n_3849)));
 assign mul_34_17_n_5577 = ((mul_34_17_n_3488 & mul_34_17_n_3801) | ((mul_34_17_n_3488 & mul_34_17_n_3489)
    | (mul_34_17_n_3489 & mul_34_17_n_3801)));
 assign mul_34_17_n_5576 = ((mul_34_17_n_3483 & mul_34_17_n_3799) | ((mul_34_17_n_3483 & mul_34_17_n_2826)
    | (mul_34_17_n_2826 & mul_34_17_n_3799)));
 assign mul_34_17_n_5575 = ((mul_34_17_n_3478 & mul_34_17_n_3798) | ((mul_34_17_n_3478 & mul_34_17_n_3479)
    | (mul_34_17_n_3479 & mul_34_17_n_3798)));
 assign mul_34_17_n_5573 = ((mul_34_17_n_3471 & mul_34_17_n_3794) | ((mul_34_17_n_3471 & mul_34_17_n_3475)
    | (mul_34_17_n_3475 & mul_34_17_n_3794)));
 assign mul_34_17_n_5572 = ((mul_34_17_n_3084 & mul_34_17_n_3665) | ((mul_34_17_n_3084 & mul_34_17_n_3085)
    | (mul_34_17_n_3085 & mul_34_17_n_3665)));
 assign mul_34_17_n_5571 = ((mul_34_17_n_3468 & mul_34_17_n_3795) | ((mul_34_17_n_3468 & mul_34_17_n_3469)
    | (mul_34_17_n_3469 & mul_34_17_n_3795)));
 assign mul_34_17_n_5570 = ((mul_34_17_n_3463 & mul_34_17_n_3793) | ((mul_34_17_n_3463 & mul_34_17_n_3464)
    | (mul_34_17_n_3464 & mul_34_17_n_3793)));
 assign mul_34_17_n_5569 = ((mul_34_17_n_4082 & mul_34_17_n_4593) | ((mul_34_17_n_4082 & mul_34_17_n_4139)
    | (mul_34_17_n_4139 & mul_34_17_n_4593)));
 assign mul_34_17_n_5568 = ((mul_34_17_n_3452 & mul_34_17_n_3789) | ((mul_34_17_n_3452 & mul_34_17_n_3453)
    | (mul_34_17_n_3453 & mul_34_17_n_3789)));
 assign mul_34_17_n_5567 = ((mul_34_17_n_3472 & mul_34_17_n_3785) | ((mul_34_17_n_3472 & mul_34_17_n_3477)
    | (mul_34_17_n_3477 & mul_34_17_n_3785)));
 assign mul_34_17_n_5566 = ((mul_34_17_n_3429 & mul_34_17_n_3782) | ((mul_34_17_n_3429 & mul_34_17_n_3438)
    | (mul_34_17_n_3438 & mul_34_17_n_3782)));
 assign mul_34_17_n_5565 = ((mul_34_17_n_3434 & mul_34_17_n_3784) | ((mul_34_17_n_3434 & mul_34_17_n_3436)
    | (mul_34_17_n_3436 & mul_34_17_n_3784)));
 assign mul_34_17_n_5564 = ((mul_34_17_n_3417 & mul_34_17_n_3771) | ((mul_34_17_n_3417 & mul_34_17_n_3419)
    | (mul_34_17_n_3419 & mul_34_17_n_3771)));
 assign mul_34_17_n_5563 = ((mul_34_17_n_3435 & mul_34_17_n_3783) | ((mul_34_17_n_3435 & mul_34_17_n_3439)
    | (mul_34_17_n_3439 & mul_34_17_n_3783)));
 assign mul_34_17_n_5562 = ((mul_34_17_n_3422 & mul_34_17_n_3779) | ((mul_34_17_n_3422 & mul_34_17_n_3424)
    | (mul_34_17_n_3424 & mul_34_17_n_3779)));
 assign mul_34_17_n_5561 = ((mul_34_17_n_3110 & mul_34_17_n_3668) | ((mul_34_17_n_3110 & mul_34_17_n_3114)
    | (mul_34_17_n_3114 & mul_34_17_n_3668)));
 assign mul_34_17_n_5559 = ((mul_34_17_n_3407 & mul_34_17_n_3878) | ((mul_34_17_n_3407 & mul_34_17_n_4529)
    | (mul_34_17_n_4529 & mul_34_17_n_3878)));
 assign mul_34_17_n_5558 = ((mul_34_17_n_3482 & mul_34_17_n_3718) | ((mul_34_17_n_3482 & mul_34_17_n_3541)
    | (mul_34_17_n_3541 & mul_34_17_n_3718)));
 assign mul_34_17_n_5557 = ((mul_34_17_n_3388 & mul_34_17_n_3770) | ((mul_34_17_n_3388 & mul_34_17_n_3390)
    | (mul_34_17_n_3390 & mul_34_17_n_3770)));
 assign mul_34_17_n_5556 = ((mul_34_17_n_3383 & mul_34_17_n_3769) | ((mul_34_17_n_3383 & mul_34_17_n_3384)
    | (mul_34_17_n_3384 & mul_34_17_n_3769)));
 assign mul_34_17_n_5555 = ((mul_34_17_n_4504 & mul_34_17_n_4655) | ((mul_34_17_n_4504 & mul_34_17_n_4508)
    | (mul_34_17_n_4508 & mul_34_17_n_4655)));
 assign mul_34_17_n_5554 = ((mul_34_17_n_3345 & mul_34_17_n_3747) | ((mul_34_17_n_3345 & mul_34_17_n_3254)
    | (mul_34_17_n_3254 & mul_34_17_n_3747)));
 assign mul_34_17_n_5553 = ((mul_34_17_n_3636 & mul_34_17_n_3680) | ((mul_34_17_n_3636 & mul_34_17_n_4135)
    | (mul_34_17_n_4135 & mul_34_17_n_3680)));
 assign mul_34_17_n_5552 = ((mul_34_17_n_4327 & mul_34_17_n_3702) | ((mul_34_17_n_4327 & mul_34_17_n_3190)
    | (mul_34_17_n_3190 & mul_34_17_n_3702)));
 assign mul_34_17_n_5551 = ((mul_34_17_n_3961 & mul_34_17_n_4727) | ((mul_34_17_n_3961 & mul_34_17_n_3639)
    | (mul_34_17_n_3639 & mul_34_17_n_4727)));
 assign mul_34_17_n_5550 = ((mul_34_17_n_4054 & mul_34_17_n_3706) | ((mul_34_17_n_4054 & mul_34_17_n_4410)
    | (mul_34_17_n_4410 & mul_34_17_n_3706)));
 assign mul_34_17_n_5549 = ((mul_34_17_n_3157 & mul_34_17_n_3684) | ((mul_34_17_n_3157 & mul_34_17_n_2838)
    | (mul_34_17_n_2838 & mul_34_17_n_3684)));
 assign mul_34_17_n_5548 = ((mul_34_17_n_3214 & mul_34_17_n_3709) | ((mul_34_17_n_3214 & mul_34_17_n_3216)
    | (mul_34_17_n_3216 & mul_34_17_n_3709)));
 assign mul_34_17_n_5547 = ((mul_34_17_n_3177 & mul_34_17_n_3700) | ((mul_34_17_n_3177 & mul_34_17_n_3184)
    | (mul_34_17_n_3184 & mul_34_17_n_3700)));
 assign mul_34_17_n_5546 = ((mul_34_17_n_3359 & mul_34_17_n_3893) | ((mul_34_17_n_3359 & mul_34_17_n_3360)
    | (mul_34_17_n_3360 & mul_34_17_n_3893)));
 assign mul_34_17_n_5545 = ((mul_34_17_n_4521 & mul_34_17_n_4725) | ((mul_34_17_n_4521 & mul_34_17_n_4048)
    | (mul_34_17_n_4048 & mul_34_17_n_4725)));
 assign mul_34_17_n_5544 = ((mul_34_17_n_3515 & mul_34_17_n_3732) | ((mul_34_17_n_3515 & mul_34_17_n_3304)
    | (mul_34_17_n_3304 & mul_34_17_n_3732)));
 assign mul_34_17_n_5543 = ((mul_34_17_n_4512 & mul_34_17_n_3919) | ((mul_34_17_n_4512 & mul_34_17_n_4514)
    | (mul_34_17_n_4514 & mul_34_17_n_3919)));
 assign mul_34_17_n_5542 = ((mul_34_17_n_3277 & mul_34_17_n_3725) | ((mul_34_17_n_3277 & mul_34_17_n_3281)
    | (mul_34_17_n_3281 & mul_34_17_n_3725)));
 assign mul_34_17_n_5541 = ((mul_34_17_n_3231 & mul_34_17_n_3708) | ((mul_34_17_n_3231 & mul_34_17_n_2817)
    | (mul_34_17_n_2817 & mul_34_17_n_3708)));
 assign mul_34_17_n_5540 = ((mul_34_17_n_3574 & mul_34_17_n_3855) | ((mul_34_17_n_3574 & mul_34_17_n_3608)
    | (mul_34_17_n_3608 & mul_34_17_n_3855)));
 assign mul_34_17_n_5539 = ((mul_34_17_n_3578 & mul_34_17_n_4609) | ((mul_34_17_n_3578 & mul_34_17_n_3329)
    | (mul_34_17_n_3329 & mul_34_17_n_4609)));
 assign mul_34_17_n_5538 = ((mul_34_17_n_3225 & mul_34_17_n_3713) | ((mul_34_17_n_3225 & mul_34_17_n_3226)
    | (mul_34_17_n_3226 & mul_34_17_n_3713)));
 assign mul_34_17_n_5537 = ((mul_34_17_n_3090 & mul_34_17_n_3666) | ((mul_34_17_n_3090 & mul_34_17_n_3644)
    | (mul_34_17_n_3644 & mul_34_17_n_3666)));
 assign mul_34_17_n_5536 = ((mul_34_17_n_4502 & mul_34_17_n_4720) | ((mul_34_17_n_4502 & mul_34_17_n_4506)
    | (mul_34_17_n_4506 & mul_34_17_n_4720)));
 assign mul_34_17_n_5535 = ((mul_34_17_n_3211 & mul_34_17_n_4760) | ((mul_34_17_n_3211 & mul_34_17_n_3217)
    | (mul_34_17_n_3217 & mul_34_17_n_4760)));
 assign mul_34_17_n_5533 = ((mul_34_17_n_3656 & mul_34_17_n_3874) | ((mul_34_17_n_3656 & mul_34_17_n_3622)
    | (mul_34_17_n_3622 & mul_34_17_n_3874)));
 assign mul_34_17_n_5531 = ((mul_34_17_n_3649 & mul_34_17_n_4605) | ((mul_34_17_n_3649 & mul_34_17_n_3648)
    | (mul_34_17_n_3648 & mul_34_17_n_4605)));
 assign mul_34_17_n_5529 = ((mul_34_17_n_3206 & mul_34_17_n_3707) | ((mul_34_17_n_3206 & mul_34_17_n_3205)
    | (mul_34_17_n_3205 & mul_34_17_n_3707)));
 assign mul_34_17_n_5527 = ((mul_34_17_n_3078 & mul_34_17_n_3705) | ((mul_34_17_n_3078 & mul_34_17_n_3093)
    | (mul_34_17_n_3093 & mul_34_17_n_3705)));
 assign mul_34_17_n_5526 = ((mul_34_17_n_3249 & mul_34_17_n_3720) | ((mul_34_17_n_3249 & mul_34_17_n_3243)
    | (mul_34_17_n_3243 & mul_34_17_n_3720)));
 assign mul_34_17_n_5525 = ((mul_34_17_n_3188 & mul_34_17_n_3699) | ((mul_34_17_n_3188 & mul_34_17_n_2815)
    | (mul_34_17_n_2815 & mul_34_17_n_3699)));
 assign mul_34_17_n_5524 = ((mul_34_17_n_4540 & mul_34_17_n_3704) | ((mul_34_17_n_4540 & mul_34_17_n_3191)
    | (mul_34_17_n_3191 & mul_34_17_n_3704)));
 assign mul_34_17_n_5523 = ((mul_34_17_n_3179 & mul_34_17_n_3696) | ((mul_34_17_n_3179 & mul_34_17_n_3178)
    | (mul_34_17_n_3178 & mul_34_17_n_3696)));
 assign mul_34_17_n_5522 = ((mul_34_17_n_3264 & mul_34_17_n_3724) | ((mul_34_17_n_3264 & mul_34_17_n_3263)
    | (mul_34_17_n_3263 & mul_34_17_n_3724)));
 assign mul_34_17_n_5521 = ((mul_34_17_n_3571 & mul_34_17_n_3831) | ((mul_34_17_n_3571 & mul_34_17_n_2828)
    | (mul_34_17_n_2828 & mul_34_17_n_3831)));
 assign mul_34_17_n_5519 = ((mul_34_17_n_4163 & mul_34_17_n_3902) | ((mul_34_17_n_4163 & mul_34_17_n_3411)
    | (mul_34_17_n_3411 & mul_34_17_n_3902)));
 assign mul_34_17_n_5518 = ((mul_34_17_n_4295 & mul_34_17_n_4662) | ((mul_34_17_n_4295 & mul_34_17_n_2734)
    | (mul_34_17_n_2734 & mul_34_17_n_4662)));
 assign mul_34_17_n_5517 = ((mul_34_17_n_4560 & mul_34_17_n_4740) | ((mul_34_17_n_4560 & mul_34_17_n_4557)
    | (mul_34_17_n_4557 & mul_34_17_n_4740)));
 assign mul_34_17_n_5515 = ((mul_34_17_n_4528 & mul_34_17_n_4564) | ((mul_34_17_n_4528 & mul_34_17_n_4400)
    | (mul_34_17_n_4400 & mul_34_17_n_4564)));
 assign mul_34_17_n_5514 = ((mul_34_17_n_4489 & mul_34_17_n_4654) | ((mul_34_17_n_4489 & mul_34_17_n_4492)
    | (mul_34_17_n_4492 & mul_34_17_n_4654)));
 assign mul_34_17_n_5513 = ((mul_34_17_n_4252 & mul_34_17_n_4738) | ((mul_34_17_n_4252 & mul_34_17_n_4552)
    | (mul_34_17_n_4552 & mul_34_17_n_4738)));
 assign mul_34_17_n_5511 = ((mul_34_17_n_4181 & mul_34_17_n_3773) | ((mul_34_17_n_4181 & mul_34_17_n_4177)
    | (mul_34_17_n_4177 & mul_34_17_n_3773)));
 assign mul_34_17_n_5509 = ((mul_34_17_n_4562 & mul_34_17_n_4741) | ((mul_34_17_n_4562 & mul_34_17_n_4117)
    | (mul_34_17_n_4117 & mul_34_17_n_4741)));
 assign mul_34_17_n_5508 = ((mul_34_17_n_4089 & mul_34_17_n_4596) | ((mul_34_17_n_4089 & mul_34_17_n_3632)
    | (mul_34_17_n_3632 & mul_34_17_n_4596)));
 assign mul_34_17_n_5507 = ((mul_34_17_n_3607 & mul_34_17_n_3911) | ((mul_34_17_n_3607 & mul_34_17_n_3108)
    | (mul_34_17_n_3108 & mul_34_17_n_3911)));
 assign mul_34_17_n_5505 = ((mul_34_17_n_3325 & mul_34_17_n_4865) | ((mul_34_17_n_3325 & mul_34_17_n_3318)
    | (mul_34_17_n_3318 & mul_34_17_n_4865)));
 assign mul_34_17_n_5504 = ((mul_34_17_n_4097 & mul_34_17_n_4617) | ((mul_34_17_n_4097 & mul_34_17_n_4397)
    | (mul_34_17_n_4397 & mul_34_17_n_4617)));
 assign mul_34_17_n_5465 = ~mul_34_17_n_5464;
 assign mul_34_17_n_5452 = ~mul_34_17_n_5451;
 assign mul_34_17_n_5433 = ~mul_34_17_n_5432;
 assign mul_34_17_n_5424 = ~mul_34_17_n_5423;
 assign mul_34_17_n_5412 = ~mul_34_17_n_5413;
 assign mul_34_17_n_5410 = ~mul_34_17_n_5411;
 assign mul_34_17_n_5409 = ((mul_34_17_n_2976 & mul_34_17_n_2702) | (mul_34_17_n_4334 & mul_34_17_n_4244));
 assign mul_34_17_n_5408 = ~(mul_34_17_n_4317 ^ mul_34_17_n_4316);
 assign mul_34_17_n_5407 = ((mul_34_17_n_2975 & mul_34_17_n_2703) | (mul_34_17_n_4314 & mul_34_17_n_4021));
 assign mul_34_17_n_5403 = ~(mul_34_17_n_4500 ^ mul_34_17_n_2939);
 assign mul_34_17_n_5500 = ~((mul_34_17_n_2993 | mul_34_17_n_2744) & (mul_34_17_n_3151 | mul_34_17_n_3022));
 assign mul_34_17_n_5396 = (mul_34_17_n_4317 ^ mul_34_17_n_4316);
 assign mul_34_17_n_5395 = (mul_34_17_n_3881 ^ mul_34_17_n_4020);
 assign mul_34_17_n_5394 = ~(mul_34_17_n_3931 ^ mul_34_17_n_3058);
 assign mul_34_17_n_5393 = (mul_34_17_n_4564 ^ mul_34_17_n_4528);
 assign mul_34_17_n_5392 = ~(mul_34_17_n_4566 ^ mul_34_17_n_4112);
 assign mul_34_17_n_5499 = ~(mul_34_17_n_4841 ^ mul_34_17_n_2957);
 assign mul_34_17_n_5391 = (mul_34_17_n_4004 ^ mul_34_17_n_4006);
 assign mul_34_17_n_5498 = (mul_34_17_n_4568 ^ mul_34_17_n_4013);
 assign mul_34_17_n_5390 = ((mul_34_17_n_2855 & mul_34_17_n_3967) | ((mul_34_17_n_2855 & mul_34_17_n_2740)
    | (mul_34_17_n_2740 & mul_34_17_n_3967)));
 assign mul_34_17_n_5389 = (mul_34_17_n_3970 ^ mul_34_17_n_4842);
 assign mul_34_17_n_5497 = (mul_34_17_n_4025 ^ mul_34_17_n_4026);
 assign mul_34_17_n_5496 = (mul_34_17_n_3884 ^ mul_34_17_n_3287);
 assign mul_34_17_n_5388 = (mul_34_17_n_3994 ^ mul_34_17_n_3996);
 assign mul_34_17_n_5495 = (mul_34_17_n_4029 ^ mul_34_17_n_4030);
 assign mul_34_17_n_5387 = (mul_34_17_n_3888 ^ mul_34_17_n_3617);
 assign mul_34_17_n_5494 = (mul_34_17_n_3088 ^ mul_34_17_n_3303);
 assign mul_34_17_n_5386 = (mul_34_17_n_4576 ^ mul_34_17_n_4034);
 assign mul_34_17_n_5385 = (mul_34_17_n_3672 ^ mul_34_17_n_3628);
 assign mul_34_17_n_5384 = (mul_34_17_n_2729 ^ mul_34_17_n_3790);
 assign mul_34_17_n_5383 = (mul_34_17_n_3399 ^ mul_34_17_n_4293);
 assign mul_34_17_n_5382 = (mul_34_17_n_4519 ^ mul_34_17_n_3212);
 assign mul_34_17_n_5493 = (mul_34_17_n_4592 ^ mul_34_17_n_4038);
 assign mul_34_17_n_5381 = (mul_34_17_n_4465 ^ mul_34_17_n_4460);
 assign mul_34_17_n_5380 = ~(mul_34_17_n_4242 ^ mul_34_17_n_4042);
 assign mul_34_17_n_5379 = (mul_34_17_n_4315 ^ mul_34_17_n_4538);
 assign mul_34_17_n_5492 = (mul_34_17_n_4730 ^ mul_34_17_n_4527);
 assign mul_34_17_n_5378 = (mul_34_17_n_3898 ^ mul_34_17_n_3105);
 assign mul_34_17_n_5377 = (mul_34_17_n_4819 ^ mul_34_17_n_4023);
 assign mul_34_17_n_5491 = (mul_34_17_n_3757 ^ mul_34_17_n_3111);
 assign mul_34_17_n_5376 = (mul_34_17_n_4106 ^ mul_34_17_n_4235);
 assign mul_34_17_n_5490 = (mul_34_17_n_4563 ^ mul_34_17_n_4558);
 assign mul_34_17_n_5489 = ~(mul_34_17_n_4813 ^ mul_34_17_n_4076);
 assign mul_34_17_n_5375 = (mul_34_17_n_3643 ^ mul_34_17_n_3089);
 assign mul_34_17_n_5488 = (mul_34_17_n_4539 ^ mul_34_17_n_4396);
 assign mul_34_17_n_5374 = (mul_34_17_n_3113 ^ mul_34_17_n_3109);
 assign mul_34_17_n_5373 = (mul_34_17_n_3079 ^ mul_34_17_n_3322);
 assign mul_34_17_n_5487 = (mul_34_17_n_4810 ^ mul_34_17_n_4443);
 assign mul_34_17_n_5372 = (mul_34_17_n_4445 ^ mul_34_17_n_4498);
 assign mul_34_17_n_5371 = (mul_34_17_n_3606 ^ mul_34_17_n_4193);
 assign mul_34_17_n_5370 = (mul_34_17_n_3490 ^ mul_34_17_n_3373);
 assign mul_34_17_n_5486 = (mul_34_17_n_4556 ^ mul_34_17_n_3991);
 assign mul_34_17_n_5369 = (mul_34_17_n_4070 ^ mul_34_17_n_4398);
 assign mul_34_17_n_5485 = (mul_34_17_n_4393 ^ mul_34_17_n_4407);
 assign mul_34_17_n_5368 = (mul_34_17_n_4549 ^ mul_34_17_n_4273);
 assign mul_34_17_n_5367 = (mul_34_17_n_4204 ^ mul_34_17_n_4233);
 assign mul_34_17_n_5366 = (mul_34_17_n_4170 ^ mul_34_17_n_4209);
 assign mul_34_17_n_5365 = ~(mul_34_17_n_4199 ^ mul_34_17_n_4490);
 assign mul_34_17_n_5364 = (mul_34_17_n_4591 ^ mul_34_17_n_3522);
 assign mul_34_17_n_5363 = (mul_34_17_n_4798 ^ mul_34_17_n_4146);
 assign mul_34_17_n_5362 = (mul_34_17_n_2818 ^ mul_34_17_n_4098);
 assign mul_34_17_n_5361 = (mul_34_17_n_4102 ^ mul_34_17_n_4063);
 assign mul_34_17_n_5360 = (mul_34_17_n_4797 ^ mul_34_17_n_4052);
 assign mul_34_17_n_5359 = (mul_34_17_n_4545 ^ mul_34_17_n_4561);
 assign mul_34_17_n_5358 = (mul_34_17_n_4795 ^ mul_34_17_n_4373);
 assign mul_34_17_n_5357 = (mul_34_17_n_4432 ^ mul_34_17_n_4430);
 assign mul_34_17_n_5356 = (mul_34_17_n_4535 ^ mul_34_17_n_4269);
 assign mul_34_17_n_5484 = (mul_34_17_n_4517 ^ mul_34_17_n_4086);
 assign mul_34_17_n_5483 = (mul_34_17_n_4494 ^ mul_34_17_n_4496);
 assign mul_34_17_n_5355 = (mul_34_17_n_4415 ^ mul_34_17_n_4471);
 assign mul_34_17_n_5482 = (mul_34_17_n_3220 ^ mul_34_17_n_3265);
 assign mul_34_17_n_5481 = (mul_34_17_n_4229 ^ mul_34_17_n_4786);
 assign mul_34_17_n_5354 = (mul_34_17_n_4387 ^ mul_34_17_n_4385);
 assign mul_34_17_n_5353 = (mul_34_17_n_4416 ^ mul_34_17_n_4417);
 assign mul_34_17_n_5352 = (mul_34_17_n_4739 ^ mul_34_17_n_4555);
 assign mul_34_17_n_5480 = (mul_34_17_n_4525 ^ mul_34_17_n_2738);
 assign mul_34_17_n_5351 = (mul_34_17_n_3275 ^ mul_34_17_n_4253);
 assign mul_34_17_n_5350 = (mul_34_17_n_4707 ^ mul_34_17_n_4363);
 assign mul_34_17_n_5349 = (mul_34_17_n_4041 ^ mul_34_17_n_4375);
 assign mul_34_17_n_5348 = (mul_34_17_n_4413 ^ mul_34_17_n_4221);
 assign mul_34_17_n_5347 = (mul_34_17_n_3761 ^ mul_34_17_n_4394);
 assign mul_34_17_n_5346 = (mul_34_17_n_3575 ^ mul_34_17_n_3899);
 assign mul_34_17_n_5479 = (mul_34_17_n_4366 ^ mul_34_17_n_4369);
 assign mul_34_17_n_5478 = (mul_34_17_n_3870 ^ mul_34_17_n_3159);
 assign mul_34_17_n_5477 = (mul_34_17_n_4354 ^ mul_34_17_n_4356);
 assign mul_34_17_n_5345 = (mul_34_17_n_4251 ^ mul_34_17_n_4257);
 assign mul_34_17_n_5344 = (mul_34_17_n_4483 ^ mul_34_17_n_4715);
 assign mul_34_17_n_5343 = (mul_34_17_n_4214 ^ mul_34_17_n_4224);
 assign mul_34_17_n_5342 = (mul_34_17_n_3194 ^ mul_34_17_n_4190);
 assign mul_34_17_n_5341 = (mul_34_17_n_3465 ^ mul_34_17_n_4507);
 assign mul_34_17_n_5339 = (mul_34_17_n_3964 ^ mul_34_17_n_4840);
 assign mul_34_17_n_5337 = ~(mul_34_17_n_4834 ^ mul_34_17_n_4833);
 assign mul_34_17_n_5476 = (mul_34_17_n_3841 ^ mul_34_17_n_4194);
 assign mul_34_17_n_5475 = (mul_34_17_n_3600 ^ mul_34_17_n_4234);
 assign mul_34_17_n_5336 = (mul_34_17_n_4109 ^ mul_34_17_n_4754);
 assign mul_34_17_n_5335 = ~(mul_34_17_n_3954 ^ mul_34_17_n_3955);
 assign mul_34_17_n_5334 = (mul_34_17_n_4148 ^ mul_34_17_n_4751);
 assign mul_34_17_n_5474 = (mul_34_17_n_4083 ^ mul_34_17_n_4090);
 assign mul_34_17_n_5332 = ~(mul_34_17_n_3037 ^ mul_34_17_n_4835);
 assign mul_34_17_n_5331 = ~(mul_34_17_n_3938 ^ mul_34_17_n_3944);
 assign mul_34_17_n_5330 = ~(mul_34_17_n_3943 ^ mul_34_17_n_3055);
 assign mul_34_17_n_5328 = (mul_34_17_n_2735 ^ mul_34_17_n_3520);
 assign mul_34_17_n_5473 = (mul_34_17_n_3993 ^ mul_34_17_n_4263);
 assign mul_34_17_n_5327 = (mul_34_17_n_3054 ^ mul_34_17_n_4099);
 assign mul_34_17_n_5472 = (mul_34_17_n_2712 ^ mul_34_17_n_4047);
 assign mul_34_17_n_5471 = (mul_34_17_n_3665 ^ mul_34_17_n_3084);
 assign mul_34_17_n_5326 = (mul_34_17_n_4039 ^ mul_34_17_n_4746);
 assign mul_34_17_n_5325 = (mul_34_17_n_4743 ^ mul_34_17_n_4019);
 assign mul_34_17_n_5470 = (mul_34_17_n_4537 ^ mul_34_17_n_3990);
 assign mul_34_17_n_5324 = (mul_34_17_n_3705 ^ mul_34_17_n_3078);
 assign mul_34_17_n_5323 = (mul_34_17_n_4077 ^ mul_34_17_n_4626);
 assign mul_34_17_n_5322 = (mul_34_17_n_4773 ^ mul_34_17_n_3321);
 assign mul_34_17_n_5321 = (mul_34_17_n_4769 ^ mul_34_17_n_4289);
 assign mul_34_17_n_5320 = (mul_34_17_n_3588 ^ mul_34_17_n_4231);
 assign mul_34_17_n_5319 = (mul_34_17_n_4223 ^ mul_34_17_n_4215);
 assign mul_34_17_n_5318 = (mul_34_17_n_4770 ^ mul_34_17_n_4300);
 assign mul_34_17_n_5317 = (mul_34_17_n_4139 ^ mul_34_17_n_4593);
 assign mul_34_17_n_5316 = (mul_34_17_n_4757 ^ mul_34_17_n_4543);
 assign mul_34_17_n_5469 = (mul_34_17_n_4532 ^ mul_34_17_n_4534);
 assign mul_34_17_n_5315 = (mul_34_17_n_3633 ^ mul_34_17_n_3616);
 assign mul_34_17_n_5314 = (mul_34_17_n_3861 ^ mul_34_17_n_2849);
 assign mul_34_17_n_5313 = (mul_34_17_n_4731 ^ mul_34_17_n_4530);
 assign mul_34_17_n_5312 = (mul_34_17_n_4341 ^ mul_34_17_n_4313);
 assign mul_34_17_n_5468 = (mul_34_17_n_2842 ^ mul_34_17_n_4584);
 assign mul_34_17_n_5311 = (mul_34_17_n_4274 ^ mul_34_17_n_4217);
 assign mul_34_17_n_5310 = (mul_34_17_n_4578 ^ mul_34_17_n_4011);
 assign mul_34_17_n_5309 = (mul_34_17_n_4414 ^ mul_34_17_n_4010);
 assign mul_34_17_n_5308 = (mul_34_17_n_4033 ^ mul_34_17_n_4028);
 assign mul_34_17_n_5307 = (mul_34_17_n_3758 ^ mul_34_17_n_4186);
 assign mul_34_17_n_5467 = (mul_34_17_n_4469 ^ mul_34_17_n_4475);
 assign mul_34_17_n_5306 = (mul_34_17_n_4737 ^ mul_34_17_n_4546);
 assign mul_34_17_n_5305 = (mul_34_17_n_4557 ^ mul_34_17_n_4560);
 assign mul_34_17_n_5466 = (mul_34_17_n_4450 ^ mul_34_17_n_4452);
 assign mul_34_17_n_5304 = (mul_34_17_n_3147 ^ mul_34_17_n_4258);
 assign mul_34_17_n_5303 = (mul_34_17_n_4062 ^ mul_34_17_n_4247);
 assign mul_34_17_n_5302 = (mul_34_17_n_4712 ^ mul_34_17_n_4481);
 assign mul_34_17_n_5301 = (mul_34_17_n_4493 ^ mul_34_17_n_4491);
 assign mul_34_17_n_5464 = ~(mul_34_17_n_4868 & mul_34_17_n_2945);
 assign mul_34_17_n_5300 = (mul_34_17_n_3145 ^ mul_34_17_n_3341);
 assign mul_34_17_n_5299 = (mul_34_17_n_3812 ^ mul_34_17_n_3507);
 assign mul_34_17_n_5298 = (mul_34_17_n_4536 ^ mul_34_17_n_3371);
 assign mul_34_17_n_5297 = ~(mul_34_17_n_3579 ^ mul_34_17_n_4422);
 assign mul_34_17_n_5296 = (mul_34_17_n_4733 ^ mul_34_17_n_4009);
 assign mul_34_17_n_5295 = ~(mul_34_17_n_3999 ^ mul_34_17_n_3513);
 assign mul_34_17_n_5294 = (mul_34_17_n_4405 ^ mul_34_17_n_3558);
 assign mul_34_17_n_5293 = (mul_34_17_n_4668 ^ mul_34_17_n_3364);
 assign mul_34_17_n_5292 = (mul_34_17_n_4499 ^ mul_34_17_n_4078);
 assign mul_34_17_n_5291 = (mul_34_17_n_4513 ^ mul_34_17_n_4511);
 assign mul_34_17_n_5290 = (mul_34_17_n_3180 ^ mul_34_17_n_4286);
 assign mul_34_17_n_5463 = (mul_34_17_n_4701 ^ mul_34_17_n_3646);
 assign mul_34_17_n_5289 = (mul_34_17_n_3438 ^ mul_34_17_n_3429);
 assign mul_34_17_n_5288 = (mul_34_17_n_3638 ^ mul_34_17_n_4053);
 assign mul_34_17_n_5287 = (mul_34_17_n_3281 ^ mul_34_17_n_3277);
 assign mul_34_17_n_5286 = (mul_34_17_n_4627 ^ mul_34_17_n_4074);
 assign mul_34_17_n_5285 = (mul_34_17_n_3625 ^ mul_34_17_n_3601);
 assign mul_34_17_n_5284 = (mul_34_17_n_3118 ^ mul_34_17_n_4456);
 assign mul_34_17_n_5283 = (mul_34_17_n_4472 ^ mul_34_17_n_4449);
 assign mul_34_17_n_5282 = (mul_34_17_n_4140 ^ mul_34_17_n_4482);
 assign mul_34_17_n_5281 = (mul_34_17_n_4547 ^ mul_34_17_n_4559);
 assign mul_34_17_n_5280 = (mul_34_17_n_4364 ^ mul_34_17_n_4365);
 assign mul_34_17_n_5279 = (mul_34_17_n_4596 ^ mul_34_17_n_3632);
 assign mul_34_17_n_5278 = (mul_34_17_n_4392 ^ mul_34_17_n_4362);
 assign mul_34_17_n_5462 = (mul_34_17_n_3127 ^ mul_34_17_n_3858);
 assign mul_34_17_n_5277 = (mul_34_17_n_4059 ^ mul_34_17_n_4292);
 assign mul_34_17_n_5461 = (mul_34_17_n_4359 ^ mul_34_17_n_4360);
 assign mul_34_17_n_5276 = (mul_34_17_n_4353 ^ mul_34_17_n_3332);
 assign mul_34_17_n_5275 = (mul_34_17_n_4583 ^ mul_34_17_n_4352);
 assign mul_34_17_n_5274 = (mul_34_17_n_4346 ^ mul_34_17_n_4672);
 assign mul_34_17_n_5273 = (mul_34_17_n_4340 ^ mul_34_17_n_4670);
 assign mul_34_17_n_5272 = (mul_34_17_n_4616 ^ mul_34_17_n_4096);
 assign mul_34_17_n_5271 = (mul_34_17_n_3106 ^ mul_34_17_n_3618);
 assign mul_34_17_n_5270 = (mul_34_17_n_4328 ^ mul_34_17_n_3653);
 assign mul_34_17_n_5269 = (mul_34_17_n_3711 ^ mul_34_17_n_3232);
 assign mul_34_17_n_5268 = (mul_34_17_n_4057 ^ mul_34_17_n_4325);
 assign mul_34_17_n_5267 = (mul_34_17_n_4615 ^ mul_34_17_n_3286);
 assign mul_34_17_n_5266 = (mul_34_17_n_4673 ^ mul_34_17_n_4320);
 assign mul_34_17_n_5265 = (mul_34_17_n_4622 ^ mul_34_17_n_4455);
 assign mul_34_17_n_5264 = (mul_34_17_n_3595 ^ mul_34_17_n_4067);
 assign mul_34_17_n_5263 = ~(mul_34_17_n_4303 ^ mul_34_17_n_4305);
 assign mul_34_17_n_5460 = (mul_34_17_n_4298 ^ mul_34_17_n_3484);
 assign mul_34_17_n_5459 = (mul_34_17_n_4296 ^ mul_34_17_n_4297);
 assign mul_34_17_n_5262 = (mul_34_17_n_4669 ^ mul_34_17_n_3992);
 assign mul_34_17_n_5261 = (mul_34_17_n_4562 ^ mul_34_17_n_4741);
 assign mul_34_17_n_5260 = (mul_34_17_n_4184 ^ mul_34_17_n_3402);
 assign mul_34_17_n_5259 = ~(mul_34_17_n_4484 ^ mul_34_17_n_2847);
 assign mul_34_17_n_5258 = (mul_34_17_n_4492 ^ mul_34_17_n_4654);
 assign mul_34_17_n_5257 = (mul_34_17_n_3842 ^ mul_34_17_n_3280);
 assign mul_34_17_n_5256 = (mul_34_17_n_3460 ^ mul_34_17_n_3458);
 assign mul_34_17_n_5255 = (mul_34_17_n_3747 ^ mul_34_17_n_3345);
 assign mul_34_17_n_5254 = (mul_34_17_n_3844 ^ mul_34_17_n_3401);
 assign mul_34_17_n_5253 = (mul_34_17_n_4036 ^ mul_34_17_n_4588);
 assign mul_34_17_n_5252 = (mul_34_17_n_4383 ^ mul_34_17_n_4380);
 assign mul_34_17_n_5251 = (mul_34_17_n_4505 ^ mul_34_17_n_4501);
 assign mul_34_17_n_5250 = (mul_34_17_n_4358 ^ mul_34_17_n_4355);
 assign mul_34_17_n_5249 = (mul_34_17_n_3573 ^ mul_34_17_n_3586);
 assign mul_34_17_n_5248 = (mul_34_17_n_4645 ^ mul_34_17_n_3294);
 assign mul_34_17_n_5247 = (mul_34_17_n_3868 ^ mul_34_17_n_3564);
 assign mul_34_17_n_5246 = (mul_34_17_n_4250 ^ mul_34_17_n_4241);
 assign mul_34_17_n_5245 = (mul_34_17_n_4641 ^ mul_34_17_n_4222);
 assign mul_34_17_n_5244 = (mul_34_17_n_4213 ^ mul_34_17_n_4639);
 assign mul_34_17_n_5243 = (mul_34_17_n_4195 ^ mul_34_17_n_3451);
 assign mul_34_17_n_5242 = (mul_34_17_n_4205 ^ mul_34_17_n_4206);
 assign mul_34_17_n_5241 = (mul_34_17_n_4084 ^ mul_34_17_n_4103);
 assign mul_34_17_n_5240 = (mul_34_17_n_4634 ^ mul_34_17_n_4196);
 assign mul_34_17_n_5239 = ~(mul_34_17_n_4457 ^ mul_34_17_n_4487);
 assign mul_34_17_n_5238 = (mul_34_17_n_4633 ^ mul_34_17_n_3441);
 assign mul_34_17_n_5237 = ~(mul_34_17_n_4277 ^ mul_34_17_n_4237);
 assign mul_34_17_n_5236 = (mul_34_17_n_3836 ^ mul_34_17_n_3548);
 assign mul_34_17_n_5235 = (mul_34_17_n_4631 ^ mul_34_17_n_3645);
 assign mul_34_17_n_5234 = (mul_34_17_n_4183 ^ mul_34_17_n_3876);
 assign mul_34_17_n_5458 = (mul_34_17_n_4611 ^ mul_34_17_n_4127);
 assign mul_34_17_n_5233 = (mul_34_17_n_4629 ^ mul_34_17_n_4182);
 assign mul_34_17_n_5457 = (mul_34_17_n_4176 ^ mul_34_17_n_3772);
 assign mul_34_17_n_5232 = (mul_34_17_n_3894 ^ mul_34_17_n_3526);
 assign mul_34_17_n_5231 = (mul_34_17_n_4108 ^ mul_34_17_n_4658);
 assign mul_34_17_n_5230 = (mul_34_17_n_3537 ^ mul_34_17_n_3533);
 assign mul_34_17_n_5229 = (mul_34_17_n_4628 ^ mul_34_17_n_4171);
 assign mul_34_17_n_5228 = (mul_34_17_n_3521 ^ mul_34_17_n_3517);
 assign mul_34_17_n_5227 = (mul_34_17_n_4115 ^ mul_34_17_n_4111);
 assign mul_34_17_n_5226 = ~(mul_34_17_n_4179 ^ mul_34_17_n_4168);
 assign mul_34_17_n_5225 = (mul_34_17_n_3477 ^ mul_34_17_n_3472);
 assign mul_34_17_n_5456 = (mul_34_17_n_2717 ^ mul_34_17_n_3320);
 assign mul_34_17_n_5224 = (mul_34_17_n_4625 ^ mul_34_17_n_4283);
 assign mul_34_17_n_5455 = (mul_34_17_n_4056 ^ mul_34_17_n_4624);
 assign mul_34_17_n_5223 = (mul_34_17_n_4623 ^ mul_34_17_n_4156);
 assign mul_34_17_n_5454 = ~(mul_34_17_n_4275 ^ mul_34_17_n_4260);
 assign mul_34_17_n_5222 = (mul_34_17_n_4147 ^ mul_34_17_n_4218);
 assign mul_34_17_n_5221 = (mul_34_17_n_4081 ^ mul_34_17_n_4635);
 assign mul_34_17_n_5220 = (mul_34_17_n_4621 ^ mul_34_17_n_4150);
 assign mul_34_17_n_5219 = (mul_34_17_n_3257 ^ mul_34_17_n_4324);
 assign mul_34_17_n_5218 = (mul_34_17_n_3511 ^ mul_34_17_n_3510);
 assign mul_34_17_n_5217 = (mul_34_17_n_4776 ^ mul_34_17_n_4374);
 assign mul_34_17_n_5453 = (mul_34_17_n_3244 ^ mul_34_17_n_4446);
 assign mul_34_17_n_5451 = (mul_34_17_n_2939 ^ mul_34_17_n_4500);
 assign mul_34_17_n_5216 = (mul_34_17_n_3681 ^ mul_34_17_n_4144);
 assign mul_34_17_n_5215 = (mul_34_17_n_3547 ^ mul_34_17_n_4597);
 assign mul_34_17_n_5214 = (mul_34_17_n_4236 ^ mul_34_17_n_4095);
 assign mul_34_17_n_5213 = (mul_34_17_n_4129 ^ mul_34_17_n_4130);
 assign mul_34_17_n_5212 = (mul_34_17_n_3338 ^ mul_34_17_n_4612);
 assign mul_34_17_n_5211 = (mul_34_17_n_4118 ^ mul_34_17_n_4610);
 assign mul_34_17_n_5210 = (mul_34_17_n_4632 ^ mul_34_17_n_3258);
 assign mul_34_17_n_5209 = (mul_34_17_n_4113 ^ mul_34_17_n_4114);
 assign mul_34_17_n_5208 = (mul_34_17_n_3493 ^ mul_34_17_n_4542);
 assign mul_34_17_n_5207 = (mul_34_17_n_3253 ^ mul_34_17_n_3252);
 assign mul_34_17_n_5206 = (mul_34_17_n_4259 ^ mul_34_17_n_4403);
 assign mul_34_17_n_5450 = ((mul_34_17_n_2845 & mul_34_17_n_3806) | ((mul_34_17_n_2845 & mul_34_17_n_2715)
    | (mul_34_17_n_2715 & mul_34_17_n_3806)));
 assign mul_34_17_n_5449 = ~(mul_34_17_n_4824 ^ mul_34_17_n_2965);
 assign mul_34_17_n_5448 = ~(mul_34_17_n_4832 ^ mul_34_17_n_2961);
 assign mul_34_17_n_5447 = ~(mul_34_17_n_4843 ^ mul_34_17_n_2951);
 assign mul_34_17_n_5446 = ~(mul_34_17_n_4830 ^ mul_34_17_n_2962);
 assign mul_34_17_n_5445 = ~(mul_34_17_n_3936 ^ mul_34_17_n_2960);
 assign mul_34_17_n_5444 = ~(mul_34_17_n_3935 ^ mul_34_17_n_2953);
 assign mul_34_17_n_5443 = (mul_34_17_n_4839 ^ mul_34_17_n_2963);
 assign mul_34_17_n_5442 = ~(mul_34_17_n_4838 ^ mul_34_17_n_2959);
 assign mul_34_17_n_5441 = ~(mul_34_17_n_3933 ^ mul_34_17_n_2954);
 assign mul_34_17_n_5440 = ~(mul_34_17_n_3929 ^ mul_34_17_n_2968);
 assign mul_34_17_n_5439 = ~(mul_34_17_n_3928 ^ mul_34_17_n_2958);
 assign mul_34_17_n_5438 = (mul_34_17_n_4809 ^ mul_34_17_n_4230);
 assign mul_34_17_n_5437 = (mul_34_17_n_4479 ^ mul_34_17_n_4480);
 assign mul_34_17_n_5436 = (mul_34_17_n_3630 ^ mul_34_17_n_4453);
 assign mul_34_17_n_5435 = (mul_34_17_n_4423 ^ mul_34_17_n_4444);
 assign mul_34_17_n_5434 = (mul_34_17_n_3097 ^ mul_34_17_n_3101);
 assign mul_34_17_n_5432 = (mul_34_17_n_4079 ^ mul_34_17_n_4069);
 assign mul_34_17_n_5431 = (mul_34_17_n_3195 ^ mul_34_17_n_4665);
 assign mul_34_17_n_5430 = (mul_34_17_n_4092 ^ mul_34_17_n_4093);
 assign mul_34_17_n_5429 = ((mul_34_17_n_2812 & mul_34_17_n_4679) | ((mul_34_17_n_2812 & mul_34_17_n_2726)
    | (mul_34_17_n_2726 & mul_34_17_n_4679)));
 assign mul_34_17_n_5428 = (mul_34_17_n_3143 ^ mul_34_17_n_3141);
 assign mul_34_17_n_5427 = (mul_34_17_n_3956 ^ mul_34_17_n_3957);
 assign mul_34_17_n_5426 = (mul_34_17_n_4270 ^ mul_34_17_n_3819);
 assign mul_34_17_n_5425 = ~(mul_34_17_n_3952 ^ mul_34_17_n_3743);
 assign mul_34_17_n_5423 = (mul_34_17_n_4550 ^ mul_34_17_n_4524);
 assign mul_34_17_n_5422 = (mul_34_17_n_4722 ^ mul_34_17_n_4509);
 assign mul_34_17_n_5421 = (mul_34_17_n_4046 ^ mul_34_17_n_4745);
 assign mul_34_17_n_5420 = ~(mul_34_17_n_2942 ^ mul_34_17_n_3774);
 assign mul_34_17_n_5205 = ~(mul_34_17_n_4837 ^ mul_34_17_n_4680);
 assign mul_34_17_n_5419 = (mul_34_17_n_2742 ^ mul_34_17_n_3736);
 assign mul_34_17_n_5418 = (mul_34_17_n_4122 ^ mul_34_17_n_4043);
 assign mul_34_17_n_5204 = ~(mul_34_17_n_4829 ^ mul_34_17_n_4828);
 assign mul_34_17_n_5417 = (mul_34_17_n_3041 ^ mul_34_17_n_4826);
 assign mul_34_17_n_5416 = (mul_34_17_n_3040 ^ mul_34_17_n_3939);
 assign mul_34_17_n_5415 = ~(mul_34_17_n_3061 ^ mul_34_17_n_3941);
 assign mul_34_17_n_5414 = ~(mul_34_17_n_3975 ^ mul_34_17_n_3932);
 assign mul_34_17_n_5413 = ~(mul_34_17_n_3750 ^ mul_34_17_n_3951);
 assign mul_34_17_n_5411 = ~(mul_34_17_n_4696 ^ mul_34_17_n_3048);
 assign mul_34_17_n_5135 = ~mul_34_17_n_5136;
 assign mul_34_17_n_5203 = ~((mul_34_17_n_4389 & mul_34_17_n_3025) | (mul_34_17_n_4049 & mul_34_17_n_3967));
 assign mul_34_17_n_5202 = ~(mul_34_17_n_4903 & mul_34_17_n_3004);
 assign mul_34_17_n_5101 = (mul_34_17_n_4554 ^ mul_34_17_n_4544);
 assign mul_34_17_n_5201 = (mul_34_17_n_3295 ^ mul_34_17_n_3299);
 assign mul_34_17_n_5100 = (mul_34_17_n_3752 ^ mul_34_17_n_4526);
 assign mul_34_17_n_5099 = (mul_34_17_n_3123 ^ mul_34_17_n_3348);
 assign mul_34_17_n_5098 = (mul_34_17_n_3134 ^ mul_34_17_n_3599);
 assign mul_34_17_n_5097 = (mul_34_17_n_3602 ^ mul_34_17_n_3102);
 assign mul_34_17_n_5096 = ~(mul_34_17_n_4220 ^ mul_34_17_n_4349);
 assign mul_34_17_n_5095 = (mul_34_17_n_3108 ^ mul_34_17_n_3607);
 assign mul_34_17_n_5200 = (mul_34_17_n_3433 ^ mul_34_17_n_3431);
 assign mul_34_17_n_5094 = (mul_34_17_n_3877 ^ mul_34_17_n_3641);
 assign mul_34_17_n_5093 = (mul_34_17_n_3224 ^ mul_34_17_n_4378);
 assign mul_34_17_n_5199 = (mul_34_17_n_3853 ^ mul_34_17_n_3597);
 assign mul_34_17_n_5092 = (mul_34_17_n_4704 ^ mul_34_17_n_3171);
 assign mul_34_17_n_5091 = (mul_34_17_n_3621 ^ mul_34_17_n_3169);
 assign mul_34_17_n_5090 = (mul_34_17_n_3664 ^ mul_34_17_n_3086);
 assign mul_34_17_n_5089 = (mul_34_17_n_3609 ^ mul_34_17_n_4734);
 assign mul_34_17_n_5088 = (mul_34_17_n_3567 ^ mul_34_17_n_3594);
 assign mul_34_17_n_5087 = (mul_34_17_n_3865 ^ mul_34_17_n_3536);
 assign mul_34_17_n_5086 = (mul_34_17_n_3732 ^ mul_34_17_n_3515);
 assign mul_34_17_n_5085 = (mul_34_17_n_3080 ^ mul_34_17_n_3130);
 assign mul_34_17_n_5084 = (mul_34_17_n_3365 ^ mul_34_17_n_4409);
 assign mul_34_17_n_5083 = (mul_34_17_n_3119 ^ mul_34_17_n_3328);
 assign mul_34_17_n_5198 = (mul_34_17_n_3426 ^ mul_34_17_n_3486);
 assign mul_34_17_n_5082 = (mul_34_17_n_3366 ^ mul_34_17_n_3140);
 assign mul_34_17_n_5081 = (mul_34_17_n_3375 ^ mul_34_17_n_4064);
 assign mul_34_17_n_5197 = (mul_34_17_n_4239 ^ mul_34_17_n_3311);
 assign mul_34_17_n_5080 = (mul_34_17_n_3585 ^ mul_34_17_n_3550);
 assign mul_34_17_n_5196 = (mul_34_17_n_3655 ^ mul_34_17_n_3155);
 assign mul_34_17_n_5079 = (mul_34_17_n_3096 ^ mul_34_17_n_3098);
 assign mul_34_17_n_5078 = (mul_34_17_n_3185 ^ mul_34_17_n_3175);
 assign mul_34_17_n_5077 = (mul_34_17_n_3149 ^ mul_34_17_n_3659);
 assign mul_34_17_n_5076 = (mul_34_17_n_3288 ^ mul_34_17_n_3285);
 assign mul_34_17_n_5195 = (mul_34_17_n_4382 ^ mul_34_17_n_3629);
 assign mul_34_17_n_5075 = (mul_34_17_n_3867 ^ mul_34_17_n_3623);
 assign mul_34_17_n_5074 = (mul_34_17_n_3611 ^ mul_34_17_n_3221);
 assign mul_34_17_n_5073 = (mul_34_17_n_4523 ^ mul_34_17_n_3326);
 assign mul_34_17_n_5072 = (mul_34_17_n_3492 ^ mul_34_17_n_3505);
 assign mul_34_17_n_5071 = (mul_34_17_n_3213 ^ mul_34_17_n_3192);
 assign mul_34_17_n_5070 = (mul_34_17_n_4285 ^ mul_34_17_n_3908);
 assign mul_34_17_n_5194 = (mul_34_17_n_3563 ^ mul_34_17_n_4137);
 assign mul_34_17_n_5069 = (mul_34_17_n_3271 ^ mul_34_17_n_4266);
 assign mul_34_17_n_5068 = (mul_34_17_n_3323 ^ mul_34_17_n_3829);
 assign mul_34_17_n_5067 = (mul_34_17_n_3544 ^ mul_34_17_n_3534);
 assign mul_34_17_n_5066 = (mul_34_17_n_3497 ^ mul_34_17_n_3568);
 assign mul_34_17_n_5065 = (mul_34_17_n_4508 ^ mul_34_17_n_4504);
 assign mul_34_17_n_5193 = (mul_34_17_n_4420 ^ mul_34_17_n_4418);
 assign mul_34_17_n_5192 = (mul_34_17_n_3610 ^ mul_34_17_n_4404);
 assign mul_34_17_n_5191 = (mul_34_17_n_4427 ^ mul_34_17_n_4424);
 assign mul_34_17_n_5064 = (mul_34_17_n_3647 ^ mul_34_17_n_3637);
 assign mul_34_17_n_5063 = (mul_34_17_n_3582 ^ mul_34_17_n_4037);
 assign mul_34_17_n_5062 = (mul_34_17_n_3273 ^ mul_34_17_n_3496);
 assign mul_34_17_n_5190 = (mul_34_17_n_3907 ^ mul_34_17_n_4141);
 assign mul_34_17_n_5189 = (mul_34_17_n_3103 ^ mul_34_17_n_3506);
 assign mul_34_17_n_5061 = (mul_34_17_n_3906 ^ mul_34_17_n_3107);
 assign mul_34_17_n_5060 = (mul_34_17_n_2825 ^ mul_34_17_n_3755);
 assign mul_34_17_n_5188 = (mul_34_17_n_3481 ^ mul_34_17_n_3584);
 assign mul_34_17_n_5187 = (mul_34_17_n_3368 ^ mul_34_17_n_3198);
 assign mul_34_17_n_5059 = (mul_34_17_n_2721 ^ mul_34_17_n_3455);
 assign mul_34_17_n_5058 = (mul_34_17_n_3411 ^ mul_34_17_n_4163);
 assign mul_34_17_n_5057 = (mul_34_17_n_4388 ^ mul_34_17_n_4377);
 assign mul_34_17_n_5056 = (mul_34_17_n_3082 ^ mul_34_17_n_4793);
 assign mul_34_17_n_5055 = (mul_34_17_n_3893 ^ mul_34_17_n_3359);
 assign mul_34_17_n_5054 = (mul_34_17_n_3354 ^ mul_34_17_n_3730);
 assign mul_34_17_n_5053 = (mul_34_17_n_3363 ^ mul_34_17_n_3361);
 assign mul_34_17_n_5186 = (mul_34_17_n_3346 ^ mul_34_17_n_3347);
 assign mul_34_17_n_5185 = (mul_34_17_n_3327 ^ mul_34_17_n_3619);
 assign mul_34_17_n_5052 = (mul_34_17_n_3885 ^ mul_34_17_n_3313);
 assign mul_34_17_n_5051 = (mul_34_17_n_4280 ^ mul_34_17_n_4278);
 assign mul_34_17_n_5050 = (mul_34_17_n_3370 ^ mul_34_17_n_3356);
 assign mul_34_17_n_5184 = (mul_34_17_n_3302 ^ mul_34_17_n_4402);
 assign mul_34_17_n_5049 = (mul_34_17_n_3462 ^ mul_34_17_n_3457);
 assign mul_34_17_n_5183 = (mul_34_17_n_3301 ^ mul_34_17_n_3298);
 assign mul_34_17_n_5182 = (mul_34_17_n_3447 ^ mul_34_17_n_3509);
 assign mul_34_17_n_5048 = (mul_34_17_n_4228 ^ mul_34_17_n_4376);
 assign mul_34_17_n_5047 = (mul_34_17_n_3278 ^ mul_34_17_n_3466);
 assign mul_34_17_n_5046 = (mul_34_17_n_4149 ^ mul_34_17_n_4462);
 assign mul_34_17_n_5045 = ~(mul_34_17_n_3454 ^ mul_34_17_n_4152);
 assign mul_34_17_n_5044 = (mul_34_17_n_3121 ^ mul_34_17_n_3565);
 assign mul_34_17_n_5043 = (mul_34_17_n_3262 ^ mul_34_17_n_3248);
 assign mul_34_17_n_5042 = (mul_34_17_n_4706 ^ mul_34_17_n_3218);
 assign mul_34_17_n_5041 = (mul_34_17_n_3988 ^ mul_34_17_n_4822);
 assign mul_34_17_n_5040 = (mul_34_17_n_2840 ^ mul_34_17_n_4411);
 assign mul_34_17_n_5181 = (mul_34_17_n_4050 ^ mul_34_17_n_4162);
 assign mul_34_17_n_5180 = (mul_34_17_n_4361 ^ mul_34_17_n_4357);
 assign mul_34_17_n_5179 = (mul_34_17_n_3446 ^ mul_34_17_n_3315);
 assign mul_34_17_n_5039 = ~(mul_34_17_n_3527 ^ mul_34_17_n_4136);
 assign mul_34_17_n_5038 = (mul_34_17_n_3652 ^ mul_34_17_n_3642);
 assign mul_34_17_n_5037 = (mul_34_17_n_3197 ^ mul_34_17_n_3358);
 assign mul_34_17_n_5178 = (mul_34_17_n_3219 ^ mul_34_17_n_3120);
 assign mul_34_17_n_5036 = (mul_34_17_n_3112 ^ mul_34_17_n_3117);
 assign mul_34_17_n_5177 = (mul_34_17_n_4518 ^ mul_34_17_n_4522);
 assign mul_34_17_n_5176 = (mul_34_17_n_4022 ^ mul_34_17_n_3186);
 assign mul_34_17_n_5035 = (mul_34_17_n_4284 ^ mul_34_17_n_4105);
 assign mul_34_17_n_5175 = (mul_34_17_n_3269 ^ mul_34_17_n_4458);
 assign mul_34_17_n_5034 = (mul_34_17_n_4529 ^ mul_34_17_n_3407);
 assign mul_34_17_n_5174 = (mul_34_17_n_3650 ^ mul_34_17_n_3406);
 assign mul_34_17_n_5033 = (mul_34_17_n_4386 ^ mul_34_17_n_3654);
 assign mul_34_17_n_5032 = (mul_34_17_n_3560 ^ mul_34_17_n_3381);
 assign mul_34_17_n_5031 = (mul_34_17_n_4708 ^ mul_34_17_n_3276);
 assign mul_34_17_n_5030 = (mul_34_17_n_4467 ^ mul_34_17_n_3376);
 assign mul_34_17_n_5029 = (mul_34_17_n_4211 ^ mul_34_17_n_3385);
 assign mul_34_17_n_5028 = (mul_34_17_n_3166 ^ mul_34_17_n_3397);
 assign mul_34_17_n_5173 = ~(mul_34_17_n_3657 ^ mul_34_17_n_2827);
 assign mul_34_17_n_5172 = (mul_34_17_n_3622 ^ mul_34_17_n_3656);
 assign mul_34_17_n_5027 = (mul_34_17_n_4756 ^ mul_34_17_n_4212);
 assign mul_34_17_n_5026 = (mul_34_17_n_3648 ^ mul_34_17_n_3649);
 assign mul_34_17_n_5025 = (mul_34_17_n_2720 ^ mul_34_17_n_3847);
 assign mul_34_17_n_5024 = (mul_34_17_n_4434 ^ mul_34_17_n_3330);
 assign mul_34_17_n_5171 = (mul_34_17_n_3317 ^ mul_34_17_n_3324);
 assign mul_34_17_n_5170 = (mul_34_17_n_3480 ^ mul_34_17_n_3674);
 assign mul_34_17_n_5023 = (mul_34_17_n_3661 ^ mul_34_17_n_3210);
 assign mul_34_17_n_5022 = (mul_34_17_n_4439 ^ mul_34_17_n_4437);
 assign mul_34_17_n_5021 = (mul_34_17_n_3500 ^ mul_34_17_n_3027);
 assign mul_34_17_n_5020 = ~(mul_34_17_n_3151 ^ mul_34_17_n_3042);
 assign mul_34_17_n_5169 = (mul_34_17_n_4143 ^ mul_34_17_n_4145);
 assign mul_34_17_n_5019 = (mul_34_17_n_4142 ^ mul_34_17_n_3624);
 assign mul_34_17_n_5168 = (mul_34_17_n_3658 ^ mul_34_17_n_3620);
 assign mul_34_17_n_5018 = (mul_34_17_n_3603 ^ mul_34_17_n_3612);
 assign mul_34_17_n_5017 = ~(mul_34_17_n_3626 ^ mul_34_17_n_4264);
 assign mul_34_17_n_5016 = (mul_34_17_n_4202 ^ mul_34_17_n_4646);
 assign mul_34_17_n_5015 = (mul_34_17_n_3420 ^ mul_34_17_n_4379);
 assign mul_34_17_n_5014 = (mul_34_17_n_2828 ^ mul_34_17_n_3831);
 assign mul_34_17_n_5013 = (mul_34_17_n_2736 ^ mul_34_17_n_3830);
 assign mul_34_17_n_5012 = (mul_34_17_n_4649 ^ mul_34_17_n_4335);
 assign mul_34_17_n_5011 = ~(mul_34_17_n_4044 ^ mul_34_17_n_4015);
 assign mul_34_17_n_5010 = (mul_34_17_n_3122 ^ mul_34_17_n_3126);
 assign mul_34_17_n_5167 = (mul_34_17_n_2730 ^ mul_34_17_n_4709);
 assign mul_34_17_n_5166 = (mul_34_17_n_2851 ^ mul_34_17_n_4598);
 assign mul_34_17_n_5009 = (mul_34_17_n_4272 ^ mul_34_17_n_3572);
 assign mul_34_17_n_5008 = (mul_34_17_n_3334 ^ mul_34_17_n_4683);
 assign mul_34_17_n_5007 = (mul_34_17_n_4711 ^ mul_34_17_n_4551);
 assign mul_34_17_n_5006 = (mul_34_17_n_4124 ^ mul_34_17_n_4126);
 assign mul_34_17_n_5005 = (mul_34_17_n_3556 ^ mul_34_17_n_3554);
 assign mul_34_17_n_5004 = (mul_34_17_n_3813 ^ mul_34_17_n_3440);
 assign mul_34_17_n_5003 = (mul_34_17_n_3576 ^ mul_34_17_n_3132);
 assign mul_34_17_n_5002 = (mul_34_17_n_3450 ^ mul_34_17_n_3843);
 assign mul_34_17_n_5001 = (mul_34_17_n_3816 ^ mul_34_17_n_3525);
 assign mul_34_17_n_5000 = (mul_34_17_n_4238 ^ mul_34_17_n_2836);
 assign mul_34_17_n_4999 = (mul_34_17_n_4477 ^ mul_34_17_n_4406);
 assign mul_34_17_n_4998 = (mul_34_17_n_4710 ^ mul_34_17_n_4476);
 assign mul_34_17_n_4997 = (mul_34_17_n_3753 ^ mul_34_17_n_3987);
 assign mul_34_17_n_4996 = (mul_34_17_n_3640 ^ mul_34_17_n_4291);
 assign mul_34_17_n_4995 = (mul_34_17_n_2734 ^ mul_34_17_n_4295);
 assign mul_34_17_n_4994 = (mul_34_17_n_4244 ^ mul_34_17_n_4334);
 assign mul_34_17_n_4993 = (mul_34_17_n_4021 ^ mul_34_17_n_4314);
 assign mul_34_17_n_4992 = (mul_34_17_n_4309 ^ mul_34_17_n_4307);
 assign mul_34_17_n_4991 = (mul_34_17_n_4132 ^ mul_34_17_n_4342);
 assign mul_34_17_n_4990 = (mul_34_17_n_4336 ^ mul_34_17_n_4332);
 assign mul_34_17_n_4989 = (mul_34_17_n_4191 ^ mul_34_17_n_4321);
 assign mul_34_17_n_4988 = (mul_34_17_n_4252 ^ mul_34_17_n_4738);
 assign mul_34_17_n_4987 = (mul_34_17_n_3788 ^ mul_34_17_n_3467);
 assign mul_34_17_n_4986 = (mul_34_17_n_3811 ^ mul_34_17_n_3516);
 assign mul_34_17_n_4985 = (mul_34_17_n_3456 ^ mul_34_17_n_3461);
 assign mul_34_17_n_4984 = (mul_34_17_n_4227 ^ mul_34_17_n_4085);
 assign mul_34_17_n_4983 = (mul_34_17_n_4249 ^ mul_34_17_n_3508);
 assign mul_34_17_n_4982 = (mul_34_17_n_4208 ^ mul_34_17_n_4210);
 assign mul_34_17_n_4981 = (mul_34_17_n_4197 ^ mul_34_17_n_4198);
 assign mul_34_17_n_4980 = (mul_34_17_n_3553 ^ mul_34_17_n_4219);
 assign mul_34_17_n_4979 = (mul_34_17_n_3827 ^ mul_34_17_n_3570);
 assign mul_34_17_n_4978 = (mul_34_17_n_4749 ^ mul_34_17_n_3104);
 assign mul_34_17_n_5165 = (mul_34_17_n_4281 ^ mul_34_17_n_3091);
 assign mul_34_17_n_4977 = (mul_34_17_n_3783 ^ mul_34_17_n_3435);
 assign mul_34_17_n_4976 = (mul_34_17_n_3170 ^ mul_34_17_n_3092);
 assign mul_34_17_n_4975 = (mul_34_17_n_3799 ^ mul_34_17_n_3483);
 assign mul_34_17_n_4974 = (mul_34_17_n_3608 ^ mul_34_17_n_3574);
 assign mul_34_17_n_4973 = (mul_34_17_n_3423 ^ mul_34_17_n_3775);
 assign mul_34_17_n_4972 = (mul_34_17_n_2732 ^ mul_34_17_n_3792);
 assign mul_34_17_n_4971 = (mul_34_17_n_3793 ^ mul_34_17_n_3463);
 assign mul_34_17_n_4970 = (mul_34_17_n_3789 ^ mul_34_17_n_3452);
 assign mul_34_17_n_4969 = (mul_34_17_n_3795 ^ mul_34_17_n_3469);
 assign mul_34_17_n_4968 = (mul_34_17_n_3801 ^ mul_34_17_n_3488);
 assign mul_34_17_n_4967 = (mul_34_17_n_3797 ^ mul_34_17_n_3474);
 assign mul_34_17_n_4966 = ~(mul_34_17_n_4724 ^ mul_34_17_n_4048);
 assign mul_34_17_n_4965 = ~(mul_34_17_n_3228 ^ mul_34_17_n_3336);
 assign mul_34_17_n_5164 = (mul_34_17_n_3424 ^ mul_34_17_n_3422);
 assign mul_34_17_n_5163 = (mul_34_17_n_3414 ^ mul_34_17_n_3410);
 assign mul_34_17_n_4964 = (mul_34_17_n_3748 ^ mul_34_17_n_3357);
 assign mul_34_17_n_4963 = (mul_34_17_n_3798 ^ mul_34_17_n_3479);
 assign mul_34_17_n_4962 = (mul_34_17_n_3425 ^ mul_34_17_n_3581);
 assign mul_34_17_n_5162 = (mul_34_17_n_3904 ^ mul_34_17_n_3415);
 assign mul_34_17_n_4961 = (mul_34_17_n_3378 ^ mul_34_17_n_2843);
 assign mul_34_17_n_4960 = (mul_34_17_n_3503 ^ mul_34_17_n_3501);
 assign mul_34_17_n_4959 = (mul_34_17_n_3413 ^ mul_34_17_n_3778);
 assign mul_34_17_n_4958 = (mul_34_17_n_3383 ^ mul_34_17_n_3384);
 assign mul_34_17_n_4957 = (mul_34_17_n_2725 ^ mul_34_17_n_4703);
 assign mul_34_17_n_4956 = (mul_34_17_n_3677 ^ mul_34_17_n_3432);
 assign mul_34_17_n_5161 = (mul_34_17_n_3449 ^ mul_34_17_n_3448);
 assign mul_34_17_n_5160 = (mul_34_17_n_3389 ^ mul_34_17_n_3387);
 assign mul_34_17_n_5159 = (mul_34_17_n_3379 ^ mul_34_17_n_3377);
 assign mul_34_17_n_5158 = (mul_34_17_n_3917 ^ mul_34_17_n_3259);
 assign mul_34_17_n_5157 = (mul_34_17_n_4167 ^ mul_34_17_n_3372);
 assign mul_34_17_n_4955 = (mul_34_17_n_3333 ^ mul_34_17_n_3339);
 assign mul_34_17_n_4954 = (mul_34_17_n_3395 ^ mul_34_17_n_3393);
 assign mul_34_17_n_5156 = (mul_34_17_n_3487 ^ mul_34_17_n_3485);
 assign mul_34_17_n_5155 = (mul_34_17_n_3255 ^ mul_34_17_n_3319);
 assign mul_34_17_n_5154 = (mul_34_17_n_4164 ^ mul_34_17_n_3442);
 assign mul_34_17_n_5153 = (mul_34_17_n_3386 ^ mul_34_17_n_3382);
 assign mul_34_17_n_4953 = (mul_34_17_n_3329 ^ mul_34_17_n_3578);
 assign mul_34_17_n_4952 = (mul_34_17_n_3226 ^ mul_34_17_n_3225);
 assign mul_34_17_n_4951 = (mul_34_17_n_3875 ^ mul_34_17_n_4027);
 assign mul_34_17_n_4950 = (mul_34_17_n_3740 ^ mul_34_17_n_3316);
 assign mul_34_17_n_4949 = (mul_34_17_n_3309 ^ mul_34_17_n_3314);
 assign mul_34_17_n_4948 = ~(mul_34_17_n_4463 ^ mul_34_17_n_3267);
 assign mul_34_17_n_4947 = (mul_34_17_n_2819 ^ mul_34_17_n_3737);
 assign mul_34_17_n_4946 = (mul_34_17_n_3434 ^ mul_34_17_n_3784);
 assign mul_34_17_n_4945 = (mul_34_17_n_3408 ^ mul_34_17_n_3409);
 assign mul_34_17_n_4944 = ~(mul_34_17_n_3289 ^ mul_34_17_n_3291);
 assign mul_34_17_n_4943 = (mul_34_17_n_3541 ^ mul_34_17_n_3718);
 assign mul_34_17_n_4942 = ~(mul_34_17_n_3297 ^ mul_34_17_n_4100);
 assign mul_34_17_n_4941 = (mul_34_17_n_3176 ^ mul_34_17_n_3676);
 assign mul_34_17_n_4940 = (mul_34_17_n_3274 ^ mul_34_17_n_3727);
 assign mul_34_17_n_4939 = (mul_34_17_n_3263 ^ mul_34_17_n_3264);
 assign mul_34_17_n_4938 = ~(mul_34_17_n_3592 ^ mul_34_17_n_4138);
 assign mul_34_17_n_4937 = ~(mul_34_17_n_4727 ^ mul_34_17_n_3639);
 assign mul_34_17_n_5152 = (mul_34_17_n_3308 ^ mul_34_17_n_3227);
 assign mul_34_17_n_4936 = (mul_34_17_n_2817 ^ mul_34_17_n_3708);
 assign mul_34_17_n_4935 = (mul_34_17_n_3243 ^ mul_34_17_n_3249);
 assign mul_34_17_n_4934 = (mul_34_17_n_3709 ^ mul_34_17_n_3214);
 assign mul_34_17_n_4933 = (mul_34_17_n_3215 ^ mul_34_17_n_3710);
 assign mul_34_17_n_4932 = (mul_34_17_n_3794 ^ mul_34_17_n_3475);
 assign mul_34_17_n_4931 = (mul_34_17_n_2835 ^ mul_34_17_n_3222);
 assign mul_34_17_n_4930 = (mul_34_17_n_2724 ^ mul_34_17_n_4777);
 assign mul_34_17_n_4929 = (mul_34_17_n_3205 ^ mul_34_17_n_3206);
 assign mul_34_17_n_5151 = (mul_34_17_n_3241 ^ mul_34_17_n_3239);
 assign mul_34_17_n_5150 = (mul_34_17_n_3076 ^ mul_34_17_n_3349);
 assign mul_34_17_n_4928 = (mul_34_17_n_3706 ^ mul_34_17_n_4054);
 assign mul_34_17_n_5149 = ~(mul_34_17_n_3200 ^ mul_34_17_n_3202);
 assign mul_34_17_n_5148 = (mul_34_17_n_3651 ^ mul_34_17_n_3261);
 assign mul_34_17_n_4927 = (mul_34_17_n_3191 ^ mul_34_17_n_4540);
 assign mul_34_17_n_4926 = (mul_34_17_n_3701 ^ mul_34_17_n_4326);
 assign mul_34_17_n_4925 = (mul_34_17_n_2815 ^ mul_34_17_n_3699);
 assign mul_34_17_n_4924 = (mul_34_17_n_3223 ^ mul_34_17_n_3189);
 assign mul_34_17_n_4923 = (mul_34_17_n_3419 ^ mul_34_17_n_3417);
 assign mul_34_17_n_5147 = (mul_34_17_n_2727 ^ mul_34_17_n_3698);
 assign mul_34_17_n_4922 = (mul_34_17_n_3700 ^ mul_34_17_n_3177);
 assign mul_34_17_n_5146 = (mul_34_17_n_3178 ^ mul_34_17_n_3179);
 assign mul_34_17_n_4921 = (mul_34_17_n_3204 ^ mul_34_17_n_4408);
 assign mul_34_17_n_4920 = (mul_34_17_n_2723 ^ mul_34_17_n_3230);
 assign mul_34_17_n_4919 = (mul_34_17_n_3217 ^ mul_34_17_n_3211);
 assign mul_34_17_n_4918 = (mul_34_17_n_3162 ^ mul_34_17_n_3164);
 assign mul_34_17_n_4917 = (mul_34_17_n_3687 ^ mul_34_17_n_3160);
 assign mul_34_17_n_4916 = (mul_34_17_n_3187 ^ mul_34_17_n_4331);
 assign mul_34_17_n_4915 = (mul_34_17_n_4750 ^ mul_34_17_n_4128);
 assign mul_34_17_n_4914 = (mul_34_17_n_3173 ^ mul_34_17_n_3174);
 assign mul_34_17_n_4913 = (mul_34_17_n_3684 ^ mul_34_17_n_3157);
 assign mul_34_17_n_5145 = (mul_34_17_n_3156 ^ mul_34_17_n_3251);
 assign mul_34_17_n_4912 = (mul_34_17_n_3821 ^ mul_34_17_n_3538);
 assign mul_34_17_n_4911 = (mul_34_17_n_3152 ^ mul_34_17_n_3351);
 assign mul_34_17_n_5144 = (mul_34_17_n_3682 ^ mul_34_17_n_3542);
 assign mul_34_17_n_4910 = (mul_34_17_n_4606 ^ mul_34_17_n_3310);
 assign mul_34_17_n_4909 = (mul_34_17_n_3679 ^ mul_34_17_n_3635);
 assign mul_34_17_n_4908 = (mul_34_17_n_3840 ^ mul_34_17_n_4448);
 assign mul_34_17_n_5143 = (mul_34_17_n_3135 ^ mul_34_17_n_4071);
 assign mul_34_17_n_5141 = ~(mul_34_17_n_4785 ^ mul_34_17_n_3047);
 assign mul_34_17_n_4907 = (mul_34_17_n_3660 ^ mul_34_17_n_3064);
 assign mul_34_17_n_5140 = ~(mul_34_17_n_3043 ^ mul_34_17_n_3751);
 assign mul_34_17_n_5139 = (mul_34_17_n_3284 ^ mul_34_17_n_3283);
 assign mul_34_17_n_5138 = (mul_34_17_n_3494 ^ mul_34_17_n_3802);
 assign mul_34_17_n_4906 = ~(mul_34_17_n_3934 ^ mul_34_17_n_3746);
 assign mul_34_17_n_5137 = (mul_34_17_n_3238 ^ mul_34_17_n_3825);
 assign mul_34_17_n_5136 = ~(mul_34_17_n_3045 ^ mul_34_17_n_3833);
 assign mul_34_17_n_5134 = ~(mul_34_17_n_3856 ^ mul_34_17_n_2820);
 assign mul_34_17_n_5133 = ~(mul_34_17_n_3950 ^ mul_34_17_n_4288);
 assign mul_34_17_n_5131 = ~(mul_34_17_n_3662 ^ mul_34_17_n_3403);
 assign mul_34_17_n_5130 = (mul_34_17_n_3256 ^ mul_34_17_n_3158);
 assign mul_34_17_n_5129 = (mul_34_17_n_3444 ^ mul_34_17_n_3421);
 assign mul_34_17_n_5128 = (mul_34_17_n_3340 ^ mul_34_17_n_3470);
 assign mul_34_17_n_5127 = (mul_34_17_n_4061 ^ mul_34_17_n_3335);
 assign mul_34_17_n_5126 = (mul_34_17_n_4674 ^ mul_34_17_n_3246);
 assign mul_34_17_n_4905 = ~(mul_34_17_n_3937 ^ mul_34_17_n_3815);
 assign mul_34_17_n_5125 = ~(mul_34_17_n_3172 ^ mul_34_17_n_3634);
 assign mul_34_17_n_5124 = ~(mul_34_17_n_4515 ^ mul_34_17_n_3128);
 assign mul_34_17_n_5122 = ~(mul_34_17_n_3726 ^ mul_34_17_n_3052);
 assign mul_34_17_n_5121 = (mul_34_17_n_4426 ^ mul_34_17_n_3445);
 assign mul_34_17_n_5120 = ((mul_34_17_n_2839 & mul_34_17_n_4696) | ((mul_34_17_n_2839 & mul_34_17_n_2713)
    | (mul_34_17_n_2713 & mul_34_17_n_4696)));
 assign mul_34_17_n_5119 = ~(mul_34_17_n_3044 ^ mul_34_17_n_4783);
 assign mul_34_17_n_5118 = ((mul_34_17_n_2844 & mul_34_17_n_4784) | ((mul_34_17_n_2844 & mul_34_17_n_2722)
    | (mul_34_17_n_2722 & mul_34_17_n_4784)));
 assign mul_34_17_n_5117 = ((mul_34_17_n_2831 & mul_34_17_n_4785) | ((mul_34_17_n_2831 & mul_34_17_n_2737)
    | (mul_34_17_n_2737 & mul_34_17_n_4785)));
 assign mul_34_17_n_5116 = ((mul_34_17_n_2821 & mul_34_17_n_3815) | ((mul_34_17_n_2821 & mul_34_17_n_2741)
    | (mul_34_17_n_2741 & mul_34_17_n_3815)));
 assign mul_34_17_n_5115 = ((mul_34_17_n_2848 & mul_34_17_n_3063) | ((mul_34_17_n_2848 & mul_34_17_n_2739)
    | (mul_34_17_n_2739 & mul_34_17_n_3063)));
 assign mul_34_17_n_5114 = ((mul_34_17_n_2854 & mul_34_17_n_3746) | ((mul_34_17_n_2854 & mul_34_17_n_2716)
    | (mul_34_17_n_2716 & mul_34_17_n_3746)));
 assign mul_34_17_n_5113 = ((mul_34_17_n_2824 & mul_34_17_n_3751) | ((mul_34_17_n_2824 & mul_34_17_n_2731)
    | (mul_34_17_n_2731 & mul_34_17_n_3751)));
 assign mul_34_17_n_5112 = ((mul_34_17_n_2814 & mul_34_17_n_3750) | ((mul_34_17_n_2814 & mul_34_17_n_2728)
    | (mul_34_17_n_2728 & mul_34_17_n_3750)));
 assign mul_34_17_n_5111 = ((mul_34_17_n_2822 & mul_34_17_n_3743) | ((mul_34_17_n_2822 & mul_34_17_n_2733)
    | (mul_34_17_n_2733 & mul_34_17_n_3743)));
 assign mul_34_17_n_5110 = (mul_34_17_n_4478 ^ mul_34_17_n_4473);
 assign mul_34_17_n_5109 = ((mul_34_17_n_2841 & mul_34_17_n_3726) | ((mul_34_17_n_2841 & mul_34_17_n_2714)
    | (mul_34_17_n_2714 & mul_34_17_n_3726)));
 assign mul_34_17_n_5108 = ((mul_34_17_n_2833 & mul_34_17_n_3833) | ((mul_34_17_n_2833 & mul_34_17_n_2719)
    | (mul_34_17_n_2719 & mul_34_17_n_3833)));
 assign mul_34_17_n_5107 = ~(mul_34_17_n_3050 ^ mul_34_17_n_3806);
 assign mul_34_17_n_4894 = ~mul_34_17_n_4893;
 assign mul_34_17_n_4890 = ~mul_34_17_n_4889;
 assign mul_34_17_n_4885 = ~mul_34_17_n_4886;
 assign mul_34_17_n_4904 = ~(mul_34_17_n_3151 & mul_34_17_n_3022);
 assign mul_34_17_n_4884 = ~(mul_34_17_n_3660 & mul_34_17_n_3064);
 assign mul_34_17_n_4903 = ~(mul_34_17_n_3847 & mul_34_17_n_3005);
 assign mul_34_17_n_4883 = ~(mul_34_17_n_4389 | mul_34_17_n_3025);
 assign mul_34_17_n_4882 = ~((mul_34_17_n_2999 | mul_34_17_n_2749) & (mul_34_17_n_2998 | mul_34_17_n_2754));
 assign mul_34_17_n_4881 = ~(mul_34_17_n_3002 | (mul_34_17_n_2752 | (mul_34_17_n_3003 | mul_34_17_n_2753)));
 assign mul_34_17_n_4880 = ~(mul_34_17_n_3061 & mul_34_17_n_3941);
 assign mul_34_17_n_4879 = ~((mul_34_17_n_3000 | mul_34_17_n_2750) & (mul_34_17_n_2997 | mul_34_17_n_2747));
 assign mul_34_17_n_4878 = ~(mul_34_17_n_3267 | mul_34_17_n_4463);
 assign mul_34_17_n_4877 = ~(mul_34_17_n_2996 | (mul_34_17_n_2751 | (mul_34_17_n_3001 | mul_34_17_n_2748)));
 assign mul_34_17_n_4876 = ~(mul_34_17_n_3267 & mul_34_17_n_4463);
 assign mul_34_17_n_4902 = ~(mul_34_17_n_3929 | mul_34_17_n_2968);
 assign mul_34_17_n_4901 = ~(mul_34_17_n_4832 | mul_34_17_n_2961);
 assign mul_34_17_n_4900 = ~(mul_34_17_n_3933 | mul_34_17_n_2954);
 assign mul_34_17_n_4899 = ~(mul_34_17_n_4824 | mul_34_17_n_2965);
 assign mul_34_17_n_4898 = ~(mul_34_17_n_3774 | mul_34_17_n_2942);
 assign mul_34_17_n_4897 = ~(mul_34_17_n_4500 | mul_34_17_n_2939);
 assign mul_34_17_n_4896 = ~(mul_34_17_n_3936 | mul_34_17_n_2960);
 assign mul_34_17_n_4895 = ~(mul_34_17_n_4843 | mul_34_17_n_2951);
 assign mul_34_17_n_4893 = ~(mul_34_17_n_4841 | mul_34_17_n_2957);
 assign mul_34_17_n_4892 = ~(mul_34_17_n_4838 | mul_34_17_n_2959);
 assign mul_34_17_n_4891 = ~(mul_34_17_n_3935 | mul_34_17_n_2953);
 assign mul_34_17_n_4889 = ~(mul_34_17_n_2995 & (mul_34_17_n_2746 & (mul_34_17_n_2994 & mul_34_17_n_2745)));
 assign mul_34_17_n_4888 = ~(mul_34_17_n_4839 | mul_34_17_n_2963);
 assign mul_34_17_n_4887 = ~(mul_34_17_n_4830 | mul_34_17_n_2962);
 assign mul_34_17_n_4886 = ~(mul_34_17_n_3928 | mul_34_17_n_2958);
 assign mul_34_17_n_4850 = ~mul_34_17_n_4849;
 assign mul_34_17_n_4875 = ((mul_34_17_n_2868 & mul_34_17_n_3039) | ((mul_34_17_n_2868 & mul_34_17_n_2743)
    | (mul_34_17_n_2743 & mul_34_17_n_3039)));
 assign mul_34_17_n_4874 = ((mul_34_17_n_1749 & mul_34_17_n_1846) | (mul_34_17_n_2989 & mul_34_17_n_436));
 assign mul_34_17_n_4873 = ((mul_34_17_n_1743 & mul_34_17_n_2266) | (mul_34_17_n_2987 & mul_34_17_n_432));
 assign mul_34_17_n_4872 = ((mul_34_17_n_1753 & mul_34_17_n_2524) | (mul_34_17_n_2985 & mul_34_17_n_445));
 assign mul_34_17_n_4871 = ((mul_34_17_n_691 & mul_34_17_n_724) | (mul_34_17_n_3007 & mul_34_17_n_483));
 assign mul_34_17_n_4870 = ((mul_34_17_n_1735 & mul_34_17_n_2218) | (mul_34_17_n_2986 & mul_34_17_n_478));
 assign mul_34_17_n_4869 = ((mul_34_17_n_1751 & mul_34_17_n_2388) | (mul_34_17_n_2983 & mul_34_17_n_428));
 assign mul_34_17_n_4868 = ((mul_34_17_n_1745 & mul_34_17_n_2258) | (mul_34_17_n_2988 & mul_34_17_n_437));
 assign mul_34_17_n_4867 = ((mul_34_17_n_685 & mul_34_17_n_768) | (mul_34_17_n_3009 & mul_34_17_n_480));
 assign mul_34_17_n_4866 = ((mul_34_17_n_681 & mul_34_17_n_869) | (mul_34_17_n_3010 & mul_34_17_n_515));
 assign mul_34_17_n_4865 = ((mul_34_17_n_1737 & mul_34_17_n_2618) | (mul_34_17_n_2980 & mul_34_17_n_433));
 assign mul_34_17_n_4864 = ((mul_34_17_n_1755 & mul_34_17_n_2657) | (mul_34_17_n_2979 & mul_34_17_n_435));
 assign mul_34_17_n_4863 = ((mul_34_17_n_1757 & mul_34_17_n_2658) | (mul_34_17_n_2990 & mul_34_17_n_448));
 assign mul_34_17_n_4862 = ((mul_34_17_n_655 & mul_34_17_n_1608) | (mul_34_17_n_2973 & mul_34_17_n_449));
 assign mul_34_17_n_4861 = ((mul_34_17_n_679 & mul_34_17_n_910) | (mul_34_17_n_3011 & mul_34_17_n_474));
 assign mul_34_17_n_4860 = ((mul_34_17_n_677 & mul_34_17_n_967) | (mul_34_17_n_3012 & mul_34_17_n_473));
 assign mul_34_17_n_4859 = ((mul_34_17_n_661 & mul_34_17_n_1374) | (mul_34_17_n_3020 & mul_34_17_n_457));
 assign mul_34_17_n_4858 = ((mul_34_17_n_663 & mul_34_17_n_1372) | (mul_34_17_n_3019 & mul_34_17_n_459));
 assign mul_34_17_n_4857 = ((mul_34_17_n_665 & mul_34_17_n_1263) | (mul_34_17_n_3018 & mul_34_17_n_460));
 assign mul_34_17_n_4856 = ((mul_34_17_n_667 & mul_34_17_n_1223) | (mul_34_17_n_3017 & mul_34_17_n_462));
 assign mul_34_17_n_4855 = ((mul_34_17_n_669 & mul_34_17_n_1139) | (mul_34_17_n_3016 & mul_34_17_n_465));
 assign mul_34_17_n_4854 = ((mul_34_17_n_671 & mul_34_17_n_1105) | (mul_34_17_n_3015 & mul_34_17_n_466));
 assign mul_34_17_n_4853 = ((mul_34_17_n_673 & mul_34_17_n_1029) | (mul_34_17_n_3021 & mul_34_17_n_468));
 assign mul_34_17_n_4852 = ((mul_34_17_n_675 & mul_34_17_n_986) | (mul_34_17_n_3013 & mul_34_17_n_470));
 assign mul_34_17_n_4851 = ((mul_34_17_n_1747 & mul_34_17_n_2288) | (mul_34_17_n_2984 & mul_34_17_n_430));
 assign mul_34_17_n_4849 = ((mul_34_17_n_687 & mul_34_17_n_707) | (mul_34_17_n_3008 & mul_34_17_n_481));
 assign mul_34_17_n_4848 = ((mul_34_17_n_1739 & mul_34_17_n_2344) | (mul_34_17_n_2981 & mul_34_17_n_444));
 assign mul_34_17_n_4847 = ((mul_34_17_n_1741 & mul_34_17_n_2442) | (mul_34_17_n_2982 & mul_34_17_n_434));
 assign mul_34_17_n_4846 = ((mul_34_17_n_659 & mul_34_17_n_1512) | (mul_34_17_n_3014 & mul_34_17_n_454));
 assign mul_34_17_n_4845 = ((mul_34_17_n_657 & mul_34_17_n_1521) | (mul_34_17_n_2977 & mul_34_17_n_452));
 assign mul_34_17_n_4836 = ~mul_34_17_n_4835;
 assign mul_34_17_n_4827 = ~mul_34_17_n_4826;
 assign mul_34_17_n_4823 = ~mul_34_17_n_4822;
 assign mul_34_17_n_4820 = ~mul_34_17_n_4819;
 assign mul_34_17_n_4814 = ~mul_34_17_n_4813;
 assign mul_34_17_n_4803 = ~mul_34_17_n_4802;
 assign mul_34_17_n_4800 = ~mul_34_17_n_4799;
 assign mul_34_17_n_4791 = ~mul_34_17_n_4790;
 assign mul_34_17_n_4784 = ~mul_34_17_n_4783;
 assign mul_34_17_n_4775 = ~mul_34_17_n_4774;
 assign mul_34_17_n_4771 = ~mul_34_17_n_4770;
 assign mul_34_17_n_4767 = ~mul_34_17_n_4766;
 assign mul_34_17_n_4755 = ~mul_34_17_n_4754;
 assign mul_34_17_n_4753 = ~mul_34_17_n_4752;
 assign mul_34_17_n_4736 = ~mul_34_17_n_4735;
 assign mul_34_17_n_4732 = ~mul_34_17_n_4731;
 assign mul_34_17_n_4725 = ~mul_34_17_n_4724;
 assign mul_34_17_n_4723 = ~mul_34_17_n_4722;
 assign mul_34_17_n_4717 = ~mul_34_17_n_4716;
 assign mul_34_17_n_4714 = ~mul_34_17_n_4713;
 assign mul_34_17_n_4690 = ~mul_34_17_n_4689;
 assign mul_34_17_n_4687 = ~mul_34_17_n_4686;
 assign mul_34_17_n_4680 = ~mul_34_17_n_4679;
 assign mul_34_17_n_4675 = ~mul_34_17_n_4674;
 assign mul_34_17_n_4666 = ~mul_34_17_n_4665;
 assign mul_34_17_n_4664 = ~mul_34_17_n_4663;
 assign mul_34_17_n_4647 = ~mul_34_17_n_4646;
 assign mul_34_17_n_4644 = ~mul_34_17_n_4643;
 assign mul_34_17_n_4619 = ~mul_34_17_n_4618;
 assign mul_34_17_n_4617 = ~mul_34_17_n_4616;
 assign mul_34_17_n_4604 = ~mul_34_17_n_4603;
 assign mul_34_17_n_4582 = ~mul_34_17_n_4581;
 assign mul_34_17_n_4579 = ~mul_34_17_n_4578;
 assign mul_34_17_n_4577 = ~mul_34_17_n_4576;
 assign mul_34_17_n_4574 = ~mul_34_17_n_4573;
 assign mul_34_17_n_4569 = ~mul_34_17_n_4568;
 assign mul_34_17_n_4567 = ~mul_34_17_n_4566;
 assign mul_34_17_n_4531 = ~mul_34_17_n_4530;
 assign mul_34_17_n_4521 = ~mul_34_17_n_4520;
 assign mul_34_17_n_4516 = ~mul_34_17_n_4515;
 assign mul_34_17_n_4514 = ~mul_34_17_n_4513;
 assign mul_34_17_n_4512 = ~mul_34_17_n_4511;
 assign mul_34_17_n_4510 = ~mul_34_17_n_4509;
 assign mul_34_17_n_4506 = ~mul_34_17_n_4505;
 assign mul_34_17_n_4502 = ~mul_34_17_n_4501;
 assign mul_34_17_n_4497 = ~mul_34_17_n_4496;
 assign mul_34_17_n_4495 = ~mul_34_17_n_4494;
 assign mul_34_17_n_4489 = ~mul_34_17_n_4488;
 assign mul_34_17_n_4485 = ~mul_34_17_n_4484;
 assign mul_34_17_n_4466 = ~mul_34_17_n_4465;
 assign mul_34_17_n_4464 = ~mul_34_17_n_4463;
 assign mul_34_17_n_4461 = ~mul_34_17_n_4460;
 assign mul_34_17_n_4459 = ~mul_34_17_n_4458;
 assign mul_34_17_n_4454 = ~mul_34_17_n_4453;
 assign mul_34_17_n_4447 = ~mul_34_17_n_4446;
 assign mul_34_17_n_4440 = ~mul_34_17_n_4439;
 assign mul_34_17_n_4438 = ~mul_34_17_n_4437;
 assign mul_34_17_n_4435 = ~mul_34_17_n_4434;
 assign mul_34_17_n_4433 = ~mul_34_17_n_4432;
 assign mul_34_17_n_4431 = ~mul_34_17_n_4430;
 assign mul_34_17_n_4428 = ~mul_34_17_n_4427;
 assign mul_34_17_n_4425 = ~mul_34_17_n_4424;
 assign mul_34_17_n_4421 = ~mul_34_17_n_4420;
 assign mul_34_17_n_4419 = ~mul_34_17_n_4418;
 assign mul_34_17_n_4390 = ~mul_34_17_n_4389;
 assign mul_34_17_n_4384 = ~mul_34_17_n_4383;
 assign mul_34_17_n_4381 = ~mul_34_17_n_4380;
 assign mul_34_17_n_4370 = ~mul_34_17_n_4369;
 assign mul_34_17_n_4367 = ~mul_34_17_n_4366;
 assign mul_34_17_n_4350 = ~mul_34_17_n_4349;
 assign mul_34_17_n_4343 = ~mul_34_17_n_4342;
 assign mul_34_17_n_4339 = ~mul_34_17_n_4338;
 assign mul_34_17_n_4337 = ~mul_34_17_n_4336;
 assign mul_34_17_n_4333 = ~mul_34_17_n_4332;
 assign mul_34_17_n_4330 = ~mul_34_17_n_4329;
 assign mul_34_17_n_4327 = ~mul_34_17_n_4326;
 assign mul_34_17_n_4322 = ~mul_34_17_n_4321;
 assign mul_34_17_n_4319 = ~mul_34_17_n_4318;
 assign mul_34_17_n_4311 = ~mul_34_17_n_4310;
 assign mul_34_17_n_4306 = ~mul_34_17_n_4305;
 assign mul_34_17_n_4304 = ~mul_34_17_n_4303;
 assign mul_34_17_n_4301 = ~mul_34_17_n_4300;
 assign mul_34_17_n_4294 = ~mul_34_17_n_4293;
 assign mul_34_17_n_4287 = ~mul_34_17_n_4286;
 assign mul_34_17_n_4276 = ~mul_34_17_n_4275;
 assign mul_34_17_n_4271 = ~mul_34_17_n_4270;
 assign mul_34_17_n_4267 = ~mul_34_17_n_4266;
 assign mul_34_17_n_4265 = ~mul_34_17_n_4264;
 assign mul_34_17_n_4261 = ~mul_34_17_n_4260;
 assign mul_34_17_n_4256 = ~mul_34_17_n_4255;
 assign mul_34_17_n_4246 = ~mul_34_17_n_4245;
 assign mul_34_17_n_4243 = ~mul_34_17_n_4242;
 assign mul_34_17_n_4240 = ~mul_34_17_n_4239;
 assign mul_34_17_n_4232 = ~mul_34_17_n_4231;
 assign mul_34_17_n_4203 = ~mul_34_17_n_4202;
 assign mul_34_17_n_4200 = ~mul_34_17_n_4199;
 assign mul_34_17_n_4192 = ~mul_34_17_n_4191;
 assign mul_34_17_n_4188 = ~mul_34_17_n_4187;
 assign mul_34_17_n_4180 = ~mul_34_17_n_4179;
 assign mul_34_17_n_4177 = ~mul_34_17_n_4176;
 assign mul_34_17_n_4169 = ~mul_34_17_n_4168;
 assign mul_34_17_n_4165 = ~mul_34_17_n_4164;
 assign mul_34_17_n_4153 = ~mul_34_17_n_4152;
 assign mul_34_17_n_4133 = ~mul_34_17_n_4132;
 assign mul_34_17_n_4110 = ~mul_34_17_n_4109;
 assign mul_34_17_n_4101 = ~mul_34_17_n_4100;
 assign mul_34_17_n_4097 = ~mul_34_17_n_4096;
 assign mul_34_17_n_4072 = ~mul_34_17_n_4071;
 assign mul_34_17_n_4068 = ~mul_34_17_n_4067;
 assign mul_34_17_n_4045 = ~mul_34_17_n_4044;
 assign mul_34_17_n_4035 = ~mul_34_17_n_4034;
 assign mul_34_17_n_4024 = ~mul_34_17_n_4023;
 assign mul_34_17_n_4018 = ~mul_34_17_n_4017;
 assign mul_34_17_n_4016 = ~mul_34_17_n_4015;
 assign mul_34_17_n_4014 = ~mul_34_17_n_4013;
 assign mul_34_17_n_4012 = ~mul_34_17_n_4011;
 assign mul_34_17_n_4007 = ~mul_34_17_n_4006;
 assign mul_34_17_n_4005 = ~mul_34_17_n_4004;
 assign mul_34_17_n_4000 = ~mul_34_17_n_3999;
 assign mul_34_17_n_3997 = ~mul_34_17_n_3996;
 assign mul_34_17_n_3995 = ~mul_34_17_n_3994;
 assign mul_34_17_n_3989 = ~mul_34_17_n_3988;
 assign mul_34_17_n_3985 = ~mul_34_17_n_3986;
 assign mul_34_17_n_3984 = ~mul_34_17_n_3983;
 assign mul_34_17_n_3982 = ~mul_34_17_n_3981;
 assign mul_34_17_n_3968 = ~mul_34_17_n_3969;
 assign mul_34_17_n_3965 = ~mul_34_17_n_3966;
 assign mul_34_17_n_3963 = ~mul_34_17_n_3964;
 assign mul_34_17_n_3960 = ~(mul_34_17_n_2850 ^ mul_34_17_n_2938);
 assign mul_34_17_n_3959 = ~(mul_34_17_n_2868 ^ mul_34_17_n_2743);
 assign mul_34_17_n_4844 = ~(mul_34_17_n_2829 ^ mul_34_17_n_2940);
 assign mul_34_17_n_3958 = ~(mul_34_17_n_2970 | mul_34_17_n_3038);
 assign mul_34_17_n_3957 = ((mul_34_17_n_688 | mul_34_17_n_652) & (mul_34_17_n_11528 | mul_34_17_n_1519));
 assign mul_34_17_n_3956 = ~((mul_34_17_n_685 & mul_34_17_n_635) | (mul_34_17_n_2931 & mul_34_17_n_788));
 assign mul_34_17_n_3955 = ~((mul_34_17_n_679 & mul_34_17_n_638) | (mul_34_17_n_2926 & mul_34_17_n_911));
 assign mul_34_17_n_3954 = ~((mul_34_17_n_1755 & mul_34_17_n_1700) | (mul_34_17_n_2898 & mul_34_17_n_2649));
 assign mul_34_17_n_3953 = ~((mul_34_17_n_661 & mul_34_17_n_647) | (mul_34_17_n_2908 & mul_34_17_n_1436));
 assign mul_34_17_n_3952 = (mul_34_17_n_2733 ^ mul_34_17_n_2822);
 assign mul_34_17_n_3951 = ~(mul_34_17_n_2728 ^ mul_34_17_n_2814);
 assign mul_34_17_n_4843 = ~((mul_34_17_n_1745 & mul_34_17_n_2481) | (mul_34_17_n_2888 & mul_34_17_n_2422));
 assign mul_34_17_n_4842 = ((mul_34_17_n_685 & mul_34_17_n_792) | (mul_34_17_n_2931 & mul_34_17_n_789));
 assign mul_34_17_n_4841 = ~((mul_34_17_n_1745 & mul_34_17_n_2340) | (mul_34_17_n_2888 & mul_34_17_n_2392));
 assign mul_34_17_n_4840 = ~((mul_34_17_n_691 & mul_34_17_n_753) | (mul_34_17_n_2936 & mul_34_17_n_699));
 assign mul_34_17_n_4839 = ((mul_34_17_n_1744 | mul_34_17_n_2161) & (mul_34_17_n_11600 | mul_34_17_n_2267));
 assign mul_34_17_n_4838 = ~((mul_34_17_n_1745 & mul_34_17_n_2119) | (mul_34_17_n_2888 & mul_34_17_n_2391));
 assign mul_34_17_n_3950 = (mul_34_17_n_2718 ^ mul_34_17_n_2832);
 assign mul_34_17_n_4837 = (mul_34_17_n_2726 ^ mul_34_17_n_2812);
 assign mul_34_17_n_4835 = ~((mul_34_17_n_1753 & mul_34_17_n_2069) | (mul_34_17_n_2878 & mul_34_17_n_1873));
 assign mul_34_17_n_4834 = ((mul_34_17_n_657 & mul_34_17_n_1520) | (mul_34_17_n_2904 & mul_34_17_n_1569));
 assign mul_34_17_n_4833 = ((mul_34_17_n_687 & mul_34_17_n_739) | (mul_34_17_n_2933 & mul_34_17_n_747));
 assign mul_34_17_n_4832 = ~((mul_34_17_n_1745 & mul_34_17_n_2115) | (mul_34_17_n_2888 & mul_34_17_n_2587));
 assign mul_34_17_n_4831 = ((mul_34_17_n_671 & mul_34_17_n_1121) | (mul_34_17_n_2918 & mul_34_17_n_1108));
 assign mul_34_17_n_4830 = ~((mul_34_17_n_1745 & mul_34_17_n_2185) | (mul_34_17_n_2888 & mul_34_17_n_2290));
 assign mul_34_17_n_3949 = ~((mul_34_17_n_671 & mul_34_17_n_642) | (mul_34_17_n_2918 & mul_34_17_n_1096));
 assign mul_34_17_n_3948 = ~((mul_34_17_n_681 & mul_34_17_n_637) | (mul_34_17_n_2928 & mul_34_17_n_854));
 assign mul_34_17_n_3947 = ~((mul_34_17_n_673 & mul_34_17_n_641) | (mul_34_17_n_2920 & mul_34_17_n_1034));
 assign mul_34_17_n_3946 = ~((mul_34_17_n_675 & mul_34_17_n_640) | (mul_34_17_n_2922 & mul_34_17_n_1010));
 assign mul_34_17_n_3945 = ~((mul_34_17_n_659 & mul_34_17_n_648) | (mul_34_17_n_2906 & mul_34_17_n_1514));
 assign mul_34_17_n_4829 = ~(mul_34_17_n_2995 & mul_34_17_n_2746);
 assign mul_34_17_n_4828 = ~(mul_34_17_n_2994 & mul_34_17_n_2745);
 assign mul_34_17_n_4826 = ~((mul_34_17_n_1755 & mul_34_17_n_2133) | (mul_34_17_n_2898 & mul_34_17_n_2588));
 assign mul_34_17_n_4825 = ~((mul_34_17_n_1737 & mul_34_17_n_2002) | (mul_34_17_n_2894 & mul_34_17_n_2627));
 assign mul_34_17_n_4824 = ~((mul_34_17_n_1745 & mul_34_17_n_2502) | (mul_34_17_n_2888 & mul_34_17_n_2682));
 assign mul_34_17_n_4822 = ((mul_34_17_n_660 | mul_34_17_n_1389) & (mul_34_17_n_11570 | mul_34_17_n_1395));
 assign mul_34_17_n_4821 = ~((mul_34_17_n_1757 & mul_34_17_n_1626) | (mul_34_17_n_2900 & mul_34_17_n_2261));
 assign mul_34_17_n_4819 = ((mul_34_17_n_670 | mul_34_17_n_1124) & (mul_34_17_n_11555 | mul_34_17_n_1094));
 assign mul_34_17_n_4818 = ~((mul_34_17_n_655 & mul_34_17_n_1641) | (mul_34_17_n_2902 & mul_34_17_n_1653));
 assign mul_34_17_n_4817 = ~((mul_34_17_n_691 & mul_34_17_n_736) | (mul_34_17_n_2936 & mul_34_17_n_738));
 assign mul_34_17_n_4816 = ~((mul_34_17_n_661 & mul_34_17_n_1410) | (mul_34_17_n_2908 & mul_34_17_n_1442));
 assign mul_34_17_n_4815 = ~((mul_34_17_n_681 & mul_34_17_n_843) | (mul_34_17_n_2928 & mul_34_17_n_874));
 assign mul_34_17_n_4813 = ((mul_34_17_n_1752 | mul_34_17_n_2201) & (mul_34_17_n_11615 | mul_34_17_n_2353));
 assign mul_34_17_n_4812 = ~((mul_34_17_n_1755 & mul_34_17_n_2219) | (mul_34_17_n_2898 & mul_34_17_n_1845));
 assign mul_34_17_n_4811 = ~((mul_34_17_n_1739 & mul_34_17_n_2159) | (mul_34_17_n_2884 & mul_34_17_n_2209));
 assign mul_34_17_n_4810 = ~((mul_34_17_n_677 & mul_34_17_n_951) | (mul_34_17_n_2924 & mul_34_17_n_954));
 assign mul_34_17_n_4809 = ~((mul_34_17_n_1755 & mul_34_17_n_2588) | (mul_34_17_n_2898 & mul_34_17_n_2676));
 assign mul_34_17_n_4808 = ((mul_34_17_n_1750 | mul_34_17_n_2437) & (mul_34_17_n_11612 | mul_34_17_n_2349));
 assign mul_34_17_n_4807 = ~((mul_34_17_n_1747 & mul_34_17_n_2647) | (mul_34_17_n_11593 & mul_34_17_n_2440));
 assign mul_34_17_n_4806 = ~((mul_34_17_n_675 & mul_34_17_n_988) | (mul_34_17_n_2922 & mul_34_17_n_1011));
 assign mul_34_17_n_4805 = ~((mul_34_17_n_661 & mul_34_17_n_1436) | (mul_34_17_n_2908 & mul_34_17_n_1437));
 assign mul_34_17_n_4804 = ~((mul_34_17_n_671 & mul_34_17_n_1118) | (mul_34_17_n_2918 & mul_34_17_n_1121));
 assign mul_34_17_n_4802 = ~((mul_34_17_n_663 & mul_34_17_n_1328) | (mul_34_17_n_2910 & mul_34_17_n_1331));
 assign mul_34_17_n_4801 = ~((mul_34_17_n_1739 & mul_34_17_n_2666) | (mul_34_17_n_2884 & mul_34_17_n_2655));
 assign mul_34_17_n_4799 = ~((mul_34_17_n_677 & mul_34_17_n_938) | (mul_34_17_n_2924 & mul_34_17_n_961));
 assign mul_34_17_n_4798 = ((mul_34_17_n_660 | mul_34_17_n_1375) & (mul_34_17_n_11570 | mul_34_17_n_1424));
 assign mul_34_17_n_4797 = ((mul_34_17_n_682 | mul_34_17_n_831) & (mul_34_17_n_11537 | mul_34_17_n_806));
 assign mul_34_17_n_4796 = ~((mul_34_17_n_1735 & mul_34_17_n_2071) | (mul_34_17_n_2896 & mul_34_17_n_2659));
 assign mul_34_17_n_4795 = ((mul_34_17_n_688 | mul_34_17_n_1519) & (mul_34_17_n_11528 | mul_34_17_n_709));
 assign mul_34_17_n_4794 = ((mul_34_17_n_657 & mul_34_17_n_1547) | (mul_34_17_n_2904 & mul_34_17_n_1525));
 assign mul_34_17_n_4793 = ((mul_34_17_n_1753 & mul_34_17_n_2567) | (mul_34_17_n_2878 & mul_34_17_n_2259));
 assign mul_34_17_n_4792 = ~((mul_34_17_n_657 & mul_34_17_n_1578) | (mul_34_17_n_2904 & mul_34_17_n_1586));
 assign mul_34_17_n_4790 = ~((mul_34_17_n_1753 & mul_34_17_n_1697) | (mul_34_17_n_2878 & mul_34_17_n_2202));
 assign mul_34_17_n_4789 = ((mul_34_17_n_1743 & mul_34_17_n_2535) | (mul_34_17_n_2882 & mul_34_17_n_2488));
 assign mul_34_17_n_4788 = ((mul_34_17_n_655 & mul_34_17_n_1639) | (mul_34_17_n_2902 & mul_34_17_n_1646));
 assign mul_34_17_n_4787 = ~((mul_34_17_n_685 & mul_34_17_n_772) | (mul_34_17_n_2931 & mul_34_17_n_771));
 assign mul_34_17_n_4786 = ((mul_34_17_n_673 & mul_34_17_n_1040) | (mul_34_17_n_2920 & mul_34_17_n_1054));
 assign mul_34_17_n_4785 = ~((mul_34_17_n_1743 & mul_34_17_n_2109) | (mul_34_17_n_2882 & mul_34_17_n_2333));
 assign mul_34_17_n_4783 = ~((mul_34_17_n_1749 & mul_34_17_n_2358) | (mul_34_17_n_2890 & mul_34_17_n_1992));
 assign mul_34_17_n_4782 = ~((mul_34_17_n_673 & mul_34_17_n_1034) | (mul_34_17_n_2920 & mul_34_17_n_1051));
 assign mul_34_17_n_4781 = ((mul_34_17_n_672 | mul_34_17_n_1015) & (mul_34_17_n_11552 | mul_34_17_n_1066));
 assign mul_34_17_n_4780 = ((mul_34_17_n_1737 & mul_34_17_n_2245) | (mul_34_17_n_2894 & mul_34_17_n_2182));
 assign mul_34_17_n_4779 = ~((mul_34_17_n_671 & mul_34_17_n_1119) | (mul_34_17_n_2918 & mul_34_17_n_1076));
 assign mul_34_17_n_4778 = ~((mul_34_17_n_675 & mul_34_17_n_995) | (mul_34_17_n_2922 & mul_34_17_n_973));
 assign mul_34_17_n_4777 = ~((mul_34_17_n_1745 & mul_34_17_n_2643) | (mul_34_17_n_2888 & mul_34_17_n_2135));
 assign mul_34_17_n_4776 = ~((mul_34_17_n_673 & mul_34_17_n_1047) | (mul_34_17_n_2920 & mul_34_17_n_1062));
 assign mul_34_17_n_4774 = ~((mul_34_17_n_663 & mul_34_17_n_1331) | (mul_34_17_n_2910 & mul_34_17_n_1350));
 assign mul_34_17_n_4773 = ~((mul_34_17_n_681 & mul_34_17_n_863) | (mul_34_17_n_2928 & mul_34_17_n_870));
 assign mul_34_17_n_4772 = ~((mul_34_17_n_673 & mul_34_17_n_1054) | (mul_34_17_n_2920 & mul_34_17_n_1060));
 assign mul_34_17_n_4770 = ((mul_34_17_n_682 | mul_34_17_n_811) & (mul_34_17_n_11537 | mul_34_17_n_815));
 assign mul_34_17_n_4769 = ~((mul_34_17_n_671 & mul_34_17_n_1095) | (mul_34_17_n_2918 & mul_34_17_n_1114));
 assign mul_34_17_n_4768 = ~((mul_34_17_n_1751 & mul_34_17_n_2580) | (mul_34_17_n_2880 & mul_34_17_n_2626));
 assign mul_34_17_n_4766 = ~((mul_34_17_n_659 & mul_34_17_n_1453) | (mul_34_17_n_2906 & mul_34_17_n_1518));
 assign mul_34_17_n_4765 = ~((mul_34_17_n_661 & mul_34_17_n_1390) | (mul_34_17_n_2908 & mul_34_17_n_1391));
 assign mul_34_17_n_4764 = ((mul_34_17_n_657 & mul_34_17_n_1588) | (mul_34_17_n_2904 & mul_34_17_n_1543));
 assign mul_34_17_n_4763 = ((mul_34_17_n_669 & mul_34_17_n_1151) | (mul_34_17_n_2916 & mul_34_17_n_1152));
 assign mul_34_17_n_4762 = ~((mul_34_17_n_687 & mul_34_17_n_749) | (mul_34_17_n_2933 & mul_34_17_n_750));
 assign mul_34_17_n_4761 = ~((mul_34_17_n_1757 & mul_34_17_n_1771) | (mul_34_17_n_2900 & mul_34_17_n_1765));
 assign mul_34_17_n_4760 = ~((mul_34_17_n_1737 & mul_34_17_n_1900) | (mul_34_17_n_2894 & mul_34_17_n_2544));
 assign mul_34_17_n_4759 = ((mul_34_17_n_688 | mul_34_17_n_696) & (mul_34_17_n_11528 | mul_34_17_n_902));
 assign mul_34_17_n_4758 = ~((mul_34_17_n_655 & mul_34_17_n_1592) | (mul_34_17_n_2902 & mul_34_17_n_1630));
 assign mul_34_17_n_4757 = ~((mul_34_17_n_681 & mul_34_17_n_858) | (mul_34_17_n_2928 & mul_34_17_n_855));
 assign mul_34_17_n_4756 = ~((mul_34_17_n_1757 & mul_34_17_n_1233) | (mul_34_17_n_2900 & mul_34_17_n_1769));
 assign mul_34_17_n_4754 = ~((mul_34_17_n_1741 & mul_34_17_n_2363) | (mul_34_17_n_2886 & mul_34_17_n_2632));
 assign mul_34_17_n_4752 = ~((mul_34_17_n_685 & mul_34_17_n_790) | (mul_34_17_n_2931 & mul_34_17_n_772));
 assign mul_34_17_n_4751 = ~((mul_34_17_n_1747 & mul_34_17_n_2426) | (mul_34_17_n_11593 & mul_34_17_n_1878));
 assign mul_34_17_n_4750 = ~((mul_34_17_n_1741 & mul_34_17_n_1853) | (mul_34_17_n_2886 & mul_34_17_n_1908));
 assign mul_34_17_n_4749 = ~((mul_34_17_n_1755 & mul_34_17_n_1889) | (mul_34_17_n_2898 & mul_34_17_n_1858));
 assign mul_34_17_n_4748 = ~((mul_34_17_n_1741 & mul_34_17_n_2406) | (mul_34_17_n_2886 & mul_34_17_n_2673));
 assign mul_34_17_n_4747 = ~((mul_34_17_n_663 & mul_34_17_n_1350) | (mul_34_17_n_2910 & mul_34_17_n_1320));
 assign mul_34_17_n_4746 = ~((mul_34_17_n_661 & mul_34_17_n_1427) | (mul_34_17_n_2908 & mul_34_17_n_1390));
 assign mul_34_17_n_4745 = ~((mul_34_17_n_665 & mul_34_17_n_1268) | (mul_34_17_n_2912 & mul_34_17_n_1299));
 assign mul_34_17_n_4744 = ~((mul_34_17_n_681 & mul_34_17_n_870) | (mul_34_17_n_2928 & mul_34_17_n_865));
 assign mul_34_17_n_4743 = ~((mul_34_17_n_679 & mul_34_17_n_885) | (mul_34_17_n_2926 & mul_34_17_n_888));
 assign mul_34_17_n_4742 = ~((mul_34_17_n_671 & mul_34_17_n_1114) | (mul_34_17_n_2918 & mul_34_17_n_1107));
 assign mul_34_17_n_4741 = ((mul_34_17_n_1734 | mul_34_17_n_2629) & (mul_34_17_n_11588 | mul_34_17_n_2601));
 assign mul_34_17_n_4740 = ((mul_34_17_n_1756 | mul_34_17_n_2096) & (mul_34_17_n_11582 | mul_34_17_n_1766));
 assign mul_34_17_n_4739 = ~((mul_34_17_n_673 & mul_34_17_n_1060) | (mul_34_17_n_2920 & mul_34_17_n_1020));
 assign mul_34_17_n_4738 = ~((mul_34_17_n_655 & mul_34_17_n_1623) | (mul_34_17_n_2902 & mul_34_17_n_1622));
 assign mul_34_17_n_4737 = ~((mul_34_17_n_691 & mul_34_17_n_738) | (mul_34_17_n_2936 & mul_34_17_n_1009));
 assign mul_34_17_n_4735 = ~((mul_34_17_n_687 & mul_34_17_n_744) | (mul_34_17_n_2933 & mul_34_17_n_695));
 assign mul_34_17_n_4734 = ~((mul_34_17_n_661 & mul_34_17_n_1426) | (mul_34_17_n_2908 & mul_34_17_n_1422));
 assign mul_34_17_n_4733 = ((mul_34_17_n_1752 | mul_34_17_n_1944) & (mul_34_17_n_11615 | mul_34_17_n_2677));
 assign mul_34_17_n_4731 = ((mul_34_17_n_668 | mul_34_17_n_1173) & (mul_34_17_n_11558 | mul_34_17_n_1134));
 assign mul_34_17_n_4730 = ((mul_34_17_n_678 | mul_34_17_n_918) & (mul_34_17_n_11543 | mul_34_17_n_896));
 assign mul_34_17_n_4729 = ~((mul_34_17_n_1745 & mul_34_17_n_2018) | (mul_34_17_n_2888 & mul_34_17_n_2651));
 assign mul_34_17_n_4728 = ~((mul_34_17_n_1737 & mul_34_17_n_2244) | (mul_34_17_n_2894 & mul_34_17_n_2697));
 assign mul_34_17_n_4727 = ((mul_34_17_n_687 & mul_34_17_n_750) | (mul_34_17_n_2933 & mul_34_17_n_743));
 assign mul_34_17_n_4726 = ~((mul_34_17_n_663 & mul_34_17_n_1366) | (mul_34_17_n_2910 & mul_34_17_n_1357));
 assign mul_34_17_n_4724 = ((mul_34_17_n_1740 | mul_34_17_n_2600) & (mul_34_17_n_11603 | mul_34_17_n_1913));
 assign mul_34_17_n_4722 = ((mul_34_17_n_1750 | mul_34_17_n_2330) & (mul_34_17_n_11612 | mul_34_17_n_2555));
 assign mul_34_17_n_4721 = ~((mul_34_17_n_1735 & mul_34_17_n_2010) | (mul_34_17_n_2896 & mul_34_17_n_2517));
 assign mul_34_17_n_4720 = ((mul_34_17_n_673 & mul_34_17_n_1020) | (mul_34_17_n_2920 & mul_34_17_n_1014));
 assign mul_34_17_n_4719 = ~((mul_34_17_n_1735 & mul_34_17_n_2602) | (mul_34_17_n_2896 & mul_34_17_n_1926));
 assign mul_34_17_n_4718 = ~((mul_34_17_n_675 & mul_34_17_n_1000) | (mul_34_17_n_2922 & mul_34_17_n_998));
 assign mul_34_17_n_4716 = ~((mul_34_17_n_679 & mul_34_17_n_881) | (mul_34_17_n_2926 & mul_34_17_n_919));
 assign mul_34_17_n_4715 = ~((mul_34_17_n_1755 & mul_34_17_n_2148) | (mul_34_17_n_2898 & mul_34_17_n_2557));
 assign mul_34_17_n_4713 = ((mul_34_17_n_1756 | mul_34_17_n_1342) & (mul_34_17_n_11582 | mul_34_17_n_1476));
 assign mul_34_17_n_4712 = ~((mul_34_17_n_679 & mul_34_17_n_905) | (mul_34_17_n_2926 & mul_34_17_n_877));
 assign mul_34_17_n_4711 = ~((mul_34_17_n_1739 & mul_34_17_n_2390) | (mul_34_17_n_2884 & mul_34_17_n_2195));
 assign mul_34_17_n_4710 = ~((mul_34_17_n_681 & mul_34_17_n_865) | (mul_34_17_n_2928 & mul_34_17_n_871));
 assign mul_34_17_n_4709 = ~((mul_34_17_n_1745 & mul_34_17_n_2149) | (mul_34_17_n_2888 & mul_34_17_n_2162));
 assign mul_34_17_n_4708 = ~((mul_34_17_n_685 & mul_34_17_n_800) | (mul_34_17_n_2931 & mul_34_17_n_767));
 assign mul_34_17_n_4707 = ~((mul_34_17_n_675 & mul_34_17_n_972) | (mul_34_17_n_2922 & mul_34_17_n_989));
 assign mul_34_17_n_4706 = ((mul_34_17_n_682 | mul_34_17_n_814) & (mul_34_17_n_11537 | mul_34_17_n_830));
 assign mul_34_17_n_4705 = ~((mul_34_17_n_1739 & mul_34_17_n_2687) | (mul_34_17_n_2884 & mul_34_17_n_2395));
 assign mul_34_17_n_4704 = ((mul_34_17_n_1736 | mul_34_17_n_2460) & (mul_34_17_n_11591 | mul_34_17_n_2332));
 assign mul_34_17_n_4703 = ~((mul_34_17_n_1745 & mul_34_17_n_2392) | (mul_34_17_n_2888 & mul_34_17_n_2361));
 assign mul_34_17_n_4702 = ((mul_34_17_n_1739 & mul_34_17_n_1955) | (mul_34_17_n_2884 & mul_34_17_n_1957));
 assign mul_34_17_n_4701 = ((mul_34_17_n_668 | mul_34_17_n_1178) & (mul_34_17_n_11558 | mul_34_17_n_1149));
 assign mul_34_17_n_4700 = ((mul_34_17_n_687 & mul_34_17_n_718) | (mul_34_17_n_2933 & mul_34_17_n_1113));
 assign mul_34_17_n_4699 = ((mul_34_17_n_663 & mul_34_17_n_1330) | (mul_34_17_n_2910 & mul_34_17_n_1322));
 assign mul_34_17_n_4698 = ~((mul_34_17_n_1739 & mul_34_17_n_2246) | (mul_34_17_n_2884 & mul_34_17_n_2309));
 assign mul_34_17_n_4697 = ((mul_34_17_n_659 & mul_34_17_n_1475) | (mul_34_17_n_2906 & mul_34_17_n_1502));
 assign mul_34_17_n_4696 = ~((mul_34_17_n_1743 & mul_34_17_n_2468) | (mul_34_17_n_2882 & mul_34_17_n_2238));
 assign mul_34_17_n_4695 = ~((mul_34_17_n_691 & mul_34_17_n_1167) | (mul_34_17_n_2936 & mul_34_17_n_754));
 assign mul_34_17_n_4694 = ~((mul_34_17_n_673 & mul_34_17_n_1019) | (mul_34_17_n_2920 & mul_34_17_n_1040));
 assign mul_34_17_n_4693 = ~((mul_34_17_n_1755 & mul_34_17_n_2557) | (mul_34_17_n_2898 & mul_34_17_n_2233));
 assign mul_34_17_n_4692 = ((mul_34_17_n_1740 | mul_34_17_n_2537) & (mul_34_17_n_11603 | mul_34_17_n_2443));
 assign mul_34_17_n_4691 = ~((mul_34_17_n_679 & mul_34_17_n_877) | (mul_34_17_n_2926 & mul_34_17_n_883));
 assign mul_34_17_n_4689 = ~((mul_34_17_n_1755 & mul_34_17_n_2385) | (mul_34_17_n_2898 & mul_34_17_n_1885));
 assign mul_34_17_n_4688 = ((mul_34_17_n_655 & mul_34_17_n_1597) | (mul_34_17_n_2902 & mul_34_17_n_1642));
 assign mul_34_17_n_4686 = ~((mul_34_17_n_691 & mul_34_17_n_734) | (mul_34_17_n_2936 & mul_34_17_n_724));
 assign mul_34_17_n_4685 = ~((mul_34_17_n_1757 & mul_34_17_n_1759) | (mul_34_17_n_2900 & mul_34_17_n_1831));
 assign mul_34_17_n_4684 = ((mul_34_17_n_682 | mul_34_17_n_825) & (mul_34_17_n_11537 | mul_34_17_n_802));
 assign mul_34_17_n_4683 = ~((mul_34_17_n_1737 & mul_34_17_n_1980) | (mul_34_17_n_2894 & mul_34_17_n_1888));
 assign mul_34_17_n_4682 = ((mul_34_17_n_682 | mul_34_17_n_808) & (mul_34_17_n_11537 | mul_34_17_n_803));
 assign mul_34_17_n_4681 = ((mul_34_17_n_1735 & mul_34_17_n_2690) | (mul_34_17_n_2896 & mul_34_17_n_2379));
 assign mul_34_17_n_4679 = ((mul_34_17_n_1742 | mul_34_17_n_2298) & (mul_34_17_n_11609 | mul_34_17_n_2489));
 assign mul_34_17_n_4678 = ~((mul_34_17_n_659 & mul_34_17_n_1479) | (mul_34_17_n_2906 & mul_34_17_n_1482));
 assign mul_34_17_n_4677 = ~((mul_34_17_n_1755 & mul_34_17_n_2014) | (mul_34_17_n_2898 & mul_34_17_n_2211));
 assign mul_34_17_n_4676 = ((mul_34_17_n_1736 | mul_34_17_n_2536) & (mul_34_17_n_11591 | mul_34_17_n_2250));
 assign mul_34_17_n_4674 = ((mul_34_17_n_1750 | mul_34_17_n_2362) & (mul_34_17_n_11612 | mul_34_17_n_2220));
 assign mul_34_17_n_4673 = ((mul_34_17_n_1749 & mul_34_17_n_2039) | (mul_34_17_n_2890 & mul_34_17_n_2272));
 assign mul_34_17_n_4672 = ((mul_34_17_n_1750 | mul_34_17_n_2526) & (mul_34_17_n_11612 | mul_34_17_n_2179));
 assign mul_34_17_n_4671 = ~((mul_34_17_n_685 & mul_34_17_n_765) | (mul_34_17_n_2931 & mul_34_17_n_762));
 assign mul_34_17_n_4670 = ((mul_34_17_n_660 | mul_34_17_n_1399) & (mul_34_17_n_11570 | mul_34_17_n_1379));
 assign mul_34_17_n_4669 = ~((mul_34_17_n_1741 & mul_34_17_n_1973) | (mul_34_17_n_2886 & mul_34_17_n_2541));
 assign mul_34_17_n_4668 = ~(mul_34_17_n_2875 ^ mul_34_17_n_2966);
 assign mul_34_17_n_4667 = ~((mul_34_17_n_669 & mul_34_17_n_1161) | (mul_34_17_n_2916 & mul_34_17_n_1166));
 assign mul_34_17_n_4665 = ((mul_34_17_n_662 | mul_34_17_n_1327) & (mul_34_17_n_11567 | mul_34_17_n_1326));
 assign mul_34_17_n_4663 = ((mul_34_17_n_1754 | mul_34_17_n_2005) & (mul_34_17_n_11585 | mul_34_17_n_2013));
 assign mul_34_17_n_4662 = ~((mul_34_17_n_1743 & mul_34_17_n_2370) | (mul_34_17_n_2882 & mul_34_17_n_2345));
 assign mul_34_17_n_4661 = ~((mul_34_17_n_671 & mul_34_17_n_1102) | (mul_34_17_n_2918 & mul_34_17_n_1117));
 assign mul_34_17_n_4660 = ~((mul_34_17_n_1735 & mul_34_17_n_2198) | (mul_34_17_n_2896 & mul_34_17_n_2417));
 assign mul_34_17_n_4659 = ((mul_34_17_n_1741 & mul_34_17_n_2616) | (mul_34_17_n_2886 & mul_34_17_n_2661));
 assign mul_34_17_n_4658 = ((mul_34_17_n_1734 | mul_34_17_n_1894) & (mul_34_17_n_11588 | mul_34_17_n_1997));
 assign mul_34_17_n_4657 = ((mul_34_17_n_1749 & mul_34_17_n_1925) | (mul_34_17_n_2890 & mul_34_17_n_2532));
 assign mul_34_17_n_4656 = ~((mul_34_17_n_681 & mul_34_17_n_853) | (mul_34_17_n_2928 & mul_34_17_n_852));
 assign mul_34_17_n_4655 = ~((mul_34_17_n_655 & mul_34_17_n_1630) | (mul_34_17_n_2902 & mul_34_17_n_1593));
 assign mul_34_17_n_4654 = ((mul_34_17_n_659 & mul_34_17_n_1509) | (mul_34_17_n_2906 & mul_34_17_n_1499));
 assign mul_34_17_n_4653 = ((mul_34_17_n_1753 & mul_34_17_n_2498) | (mul_34_17_n_2878 & mul_34_17_n_2319));
 assign mul_34_17_n_4652 = ~(mul_34_17_n_2865 ^ mul_34_17_n_2956);
 assign mul_34_17_n_4651 = ~((mul_34_17_n_691 & mul_34_17_n_721) | (mul_34_17_n_2936 & mul_34_17_n_1167));
 assign mul_34_17_n_4650 = ((mul_34_17_n_1753 & mul_34_17_n_2146) | (mul_34_17_n_2878 & mul_34_17_n_2622));
 assign mul_34_17_n_4649 = ~((mul_34_17_n_1753 & mul_34_17_n_2444) | (mul_34_17_n_2878 & mul_34_17_n_1970));
 assign mul_34_17_n_4648 = ((mul_34_17_n_1755 & mul_34_17_n_2547) | (mul_34_17_n_2898 & mul_34_17_n_2396));
 assign mul_34_17_n_4646 = ((mul_34_17_n_1754 | mul_34_17_n_1967) & (mul_34_17_n_11585 | mul_34_17_n_2090));
 assign mul_34_17_n_4645 = ~((mul_34_17_n_1757 & mul_34_17_n_1063) | (mul_34_17_n_2900 & mul_34_17_n_1233));
 assign mul_34_17_n_4643 = ~((mul_34_17_n_1747 & mul_34_17_n_2691) | (mul_34_17_n_11593 & mul_34_17_n_2366));
 assign mul_34_17_n_4642 = ((mul_34_17_n_673 & mul_34_17_n_1049) | (mul_34_17_n_2920 & mul_34_17_n_1039));
 assign mul_34_17_n_4641 = ((mul_34_17_n_1751 & mul_34_17_n_2365) | (mul_34_17_n_2880 & mul_34_17_n_2457));
 assign mul_34_17_n_4640 = ((mul_34_17_n_1751 & mul_34_17_n_2326) | (mul_34_17_n_2880 & mul_34_17_n_2459));
 assign mul_34_17_n_4639 = ((mul_34_17_n_677 & mul_34_17_n_957) | (mul_34_17_n_2924 & mul_34_17_n_943));
 assign mul_34_17_n_4638 = ((mul_34_17_n_1750 | mul_34_17_n_2224) & (mul_34_17_n_11612 | mul_34_17_n_2342));
 assign mul_34_17_n_4637 = ~((mul_34_17_n_673 & mul_34_17_n_1036) | (mul_34_17_n_2920 & mul_34_17_n_1047));
 assign mul_34_17_n_4636 = ((mul_34_17_n_1735 & mul_34_17_n_2528) | (mul_34_17_n_2896 & mul_34_17_n_2455));
 assign mul_34_17_n_4635 = ~((mul_34_17_n_1747 & mul_34_17_n_2453) | (mul_34_17_n_11593 & mul_34_17_n_2472));
 assign mul_34_17_n_4634 = ~((mul_34_17_n_663 & mul_34_17_n_1315) | (mul_34_17_n_2910 & mul_34_17_n_1354));
 assign mul_34_17_n_4633 = ~((mul_34_17_n_681 & mul_34_17_n_873) | (mul_34_17_n_2928 & mul_34_17_n_861));
 assign mul_34_17_n_4632 = ((mul_34_17_n_684 | mul_34_17_n_791) & (mul_34_17_n_11534 | mul_34_17_n_775));
 assign mul_34_17_n_4631 = ~((mul_34_17_n_661 & mul_34_17_n_1434) | (mul_34_17_n_2908 & mul_34_17_n_1419));
 assign mul_34_17_n_4630 = ((mul_34_17_n_1748 | mul_34_17_n_2237) & (mul_34_17_n_11597 | mul_34_17_n_2253));
 assign mul_34_17_n_4629 = ((mul_34_17_n_682 | mul_34_17_n_813) & (mul_34_17_n_11537 | mul_34_17_n_814));
 assign mul_34_17_n_4628 = ~((mul_34_17_n_659 & mul_34_17_n_1513) | (mul_34_17_n_2906 & mul_34_17_n_1460));
 assign mul_34_17_n_4627 = ((mul_34_17_n_1756 | mul_34_17_n_727) & (mul_34_17_n_11582 | mul_34_17_n_1678));
 assign mul_34_17_n_4626 = ((mul_34_17_n_1736 | mul_34_17_n_2376) & (mul_34_17_n_11591 | mul_34_17_n_1940));
 assign mul_34_17_n_4625 = ~((mul_34_17_n_1755 & mul_34_17_n_2452) | (mul_34_17_n_2898 & mul_34_17_n_2041));
 assign mul_34_17_n_4624 = ~((mul_34_17_n_1739 & mul_34_17_n_2564) | (mul_34_17_n_2884 & mul_34_17_n_2246));
 assign mul_34_17_n_4623 = ~((mul_34_17_n_661 & mul_34_17_n_1419) | (mul_34_17_n_2908 & mul_34_17_n_1397));
 assign mul_34_17_n_4622 = ~((mul_34_17_n_667 & mul_34_17_n_1186) | (mul_34_17_n_2914 & mul_34_17_n_1193));
 assign mul_34_17_n_4621 = ~((mul_34_17_n_675 & mul_34_17_n_983) | (mul_34_17_n_2922 & mul_34_17_n_1008));
 assign mul_34_17_n_4620 = ~((mul_34_17_n_682 | mul_34_17_n_822) & (mul_34_17_n_11537 | mul_34_17_n_805));
 assign mul_34_17_n_4618 = ~((mul_34_17_n_675 & mul_34_17_n_993) | (mul_34_17_n_2922 & mul_34_17_n_997));
 assign mul_34_17_n_4616 = ~((mul_34_17_n_655 & mul_34_17_n_1595) | (mul_34_17_n_2902 & mul_34_17_n_1658));
 assign mul_34_17_n_4615 = ~((mul_34_17_n_1749 & mul_34_17_n_1928) | (mul_34_17_n_2890 & mul_34_17_n_1925));
 assign mul_34_17_n_4614 = ~((mul_34_17_n_687 & mul_34_17_n_717) | (mul_34_17_n_2933 & mul_34_17_n_711));
 assign mul_34_17_n_4613 = ((mul_34_17_n_678 | mul_34_17_n_906) & (mul_34_17_n_11543 | mul_34_17_n_904));
 assign mul_34_17_n_4612 = ~((mul_34_17_n_1749 & mul_34_17_n_2254) | (mul_34_17_n_2890 & mul_34_17_n_2604));
 assign mul_34_17_n_4611 = ~((mul_34_17_n_673 & mul_34_17_n_1038) | (mul_34_17_n_2920 & mul_34_17_n_1019));
 assign mul_34_17_n_4610 = ~((mul_34_17_n_1735 & mul_34_17_n_2316) | (mul_34_17_n_2896 & mul_34_17_n_2071));
 assign mul_34_17_n_4609 = ~((mul_34_17_n_1739 & mul_34_17_n_2187) | (mul_34_17_n_2884 & mul_34_17_n_2339));
 assign mul_34_17_n_4608 = ~((mul_34_17_n_661 & mul_34_17_n_1425) | (mul_34_17_n_2908 & mul_34_17_n_1428));
 assign mul_34_17_n_4607 = ((mul_34_17_n_654 | mul_34_17_n_1647) & (mul_34_17_n_11579 | mul_34_17_n_1601));
 assign mul_34_17_n_4606 = ~((mul_34_17_n_1741 & mul_34_17_n_1939) | (mul_34_17_n_2886 & mul_34_17_n_2484));
 assign mul_34_17_n_4605 = ~((mul_34_17_n_1737 & mul_34_17_n_2222) | (mul_34_17_n_2894 & mul_34_17_n_2503));
 assign mul_34_17_n_4603 = ~((mul_34_17_n_659 & mul_34_17_n_1484) | (mul_34_17_n_2906 & mul_34_17_n_1492));
 assign mul_34_17_n_4602 = ~((mul_34_17_n_1745 & mul_34_17_n_2642) | (mul_34_17_n_2888 & mul_34_17_n_2545));
 assign mul_34_17_n_4601 = ~((mul_34_17_n_685 & mul_34_17_n_760) | (mul_34_17_n_2931 & mul_34_17_n_768));
 assign mul_34_17_n_4600 = ((mul_34_17_n_1750 | mul_34_17_n_1907) & (mul_34_17_n_11612 | mul_34_17_n_2675));
 assign mul_34_17_n_4599 = ~((mul_34_17_n_661 & mul_34_17_n_1421) | (mul_34_17_n_2908 & mul_34_17_n_1423));
 assign mul_34_17_n_4598 = ~((mul_34_17_n_1749 & mul_34_17_n_2341) | (mul_34_17_n_2890 & mul_34_17_n_2684));
 assign mul_34_17_n_4597 = ((mul_34_17_n_1738 | mul_34_17_n_2624) & (mul_34_17_n_11606 | mul_34_17_n_2487));
 assign mul_34_17_n_4596 = ((mul_34_17_n_690 | mul_34_17_n_719) & (mul_34_17_n_11525 | mul_34_17_n_1057));
 assign mul_34_17_n_4595 = ((mul_34_17_n_1737 & mul_34_17_n_2429) | (mul_34_17_n_2894 & mul_34_17_n_2223));
 assign mul_34_17_n_4594 = ~((mul_34_17_n_1741 & mul_34_17_n_2461) | (mul_34_17_n_2886 & mul_34_17_n_2140));
 assign mul_34_17_n_4593 = ((mul_34_17_n_1756 | mul_34_17_n_2377) & (mul_34_17_n_11582 | mul_34_17_n_727));
 assign mul_34_17_n_4592 = ((mul_34_17_n_684 | mul_34_17_n_761) & (mul_34_17_n_11534 | mul_34_17_n_759));
 assign mul_34_17_n_4591 = ~((mul_34_17_n_681 & mul_34_17_n_854) | (mul_34_17_n_2928 & mul_34_17_n_856));
 assign mul_34_17_n_4590 = ~((mul_34_17_n_1757 & mul_34_17_n_955) | (mul_34_17_n_2900 & mul_34_17_n_2615));
 assign mul_34_17_n_4589 = ((mul_34_17_n_672 | mul_34_17_n_1035) & (mul_34_17_n_11552 | mul_34_17_n_1037));
 assign mul_34_17_n_4588 = ~((mul_34_17_n_1747 & mul_34_17_n_1990) | (mul_34_17_n_11593 & mul_34_17_n_2381));
 assign mul_34_17_n_4587 = ~((mul_34_17_n_1755 & mul_34_17_n_2252) | (mul_34_17_n_2898 & mul_34_17_n_2483));
 assign mul_34_17_n_4586 = ((mul_34_17_n_660 | mul_34_17_n_1411) & (mul_34_17_n_11570 | mul_34_17_n_1412));
 assign mul_34_17_n_4585 = ~((mul_34_17_n_1741 & mul_34_17_n_1924) | (mul_34_17_n_2886 & mul_34_17_n_1989));
 assign mul_34_17_n_4584 = ((mul_34_17_n_664 | mul_34_17_n_1304) & (mul_34_17_n_11564 | mul_34_17_n_1291));
 assign mul_34_17_n_4583 = ~((mul_34_17_n_655 & mul_34_17_n_1628) | (mul_34_17_n_2902 & mul_34_17_n_1592));
 assign mul_34_17_n_4581 = ~((mul_34_17_n_1743 & mul_34_17_n_2305) | (mul_34_17_n_2882 & mul_34_17_n_2695));
 assign mul_34_17_n_4580 = ((mul_34_17_n_1745 & mul_34_17_n_2175) | (mul_34_17_n_2888 & mul_34_17_n_2165));
 assign mul_34_17_n_4578 = ((mul_34_17_n_682 | mul_34_17_n_819) & (mul_34_17_n_11537 | mul_34_17_n_813));
 assign mul_34_17_n_4576 = ((mul_34_17_n_676 | mul_34_17_n_927) & (mul_34_17_n_11546 | mul_34_17_n_964));
 assign mul_34_17_n_4575 = ~((mul_34_17_n_667 & mul_34_17_n_1244) | (mul_34_17_n_2914 & mul_34_17_n_1206));
 assign mul_34_17_n_4573 = ((mul_34_17_n_666 | mul_34_17_n_1203) & (mul_34_17_n_11561 | mul_34_17_n_1239));
 assign mul_34_17_n_4572 = ((mul_34_17_n_1734 | mul_34_17_n_2049) & (mul_34_17_n_11588 | mul_34_17_n_2031));
 assign mul_34_17_n_4571 = ~((mul_34_17_n_1745 & mul_34_17_n_1968) | (mul_34_17_n_2888 & mul_34_17_n_1920));
 assign mul_34_17_n_4570 = ~((mul_34_17_n_656 | mul_34_17_n_1534) & (mul_34_17_n_11576 | mul_34_17_n_1545));
 assign mul_34_17_n_4568 = ~((mul_34_17_n_1739 & mul_34_17_n_2328) | (mul_34_17_n_2884 & mul_34_17_n_2354));
 assign mul_34_17_n_4566 = ((mul_34_17_n_1750 | mul_34_17_n_2067) & (mul_34_17_n_11612 | mul_34_17_n_2413));
 assign mul_34_17_n_4565 = ((mul_34_17_n_1739 & mul_34_17_n_2352) | (mul_34_17_n_2884 & mul_34_17_n_2625));
 assign mul_34_17_n_4564 = ((mul_34_17_n_664 | mul_34_17_n_1296) & (mul_34_17_n_11564 | mul_34_17_n_1281));
 assign mul_34_17_n_4563 = ((mul_34_17_n_662 | mul_34_17_n_1319) & (mul_34_17_n_11567 | mul_34_17_n_1335));
 assign mul_34_17_n_4562 = ((mul_34_17_n_658 | mul_34_17_n_1517) & (mul_34_17_n_11573 | mul_34_17_n_1457));
 assign mul_34_17_n_4561 = ~((mul_34_17_n_675 & mul_34_17_n_997) | (mul_34_17_n_2922 & mul_34_17_n_995));
 assign mul_34_17_n_4560 = ((mul_34_17_n_1740 | mul_34_17_n_1695) & (mul_34_17_n_11603 | mul_34_17_n_2600));
 assign mul_34_17_n_4559 = ~((mul_34_17_n_1739 & mul_34_17_n_2655) | (mul_34_17_n_2884 & mul_34_17_n_1955));
 assign mul_34_17_n_4558 = ((mul_34_17_n_660 | mul_34_17_n_1403) & (mul_34_17_n_11570 | mul_34_17_n_1405));
 assign mul_34_17_n_4557 = ((mul_34_17_n_666 | mul_34_17_n_1194) & (mul_34_17_n_11561 | mul_34_17_n_1243));
 assign mul_34_17_n_4556 = ~((mul_34_17_n_675 & mul_34_17_n_1002) | (mul_34_17_n_2922 & mul_34_17_n_968));
 assign mul_34_17_n_4555 = ~((mul_34_17_n_663 & mul_34_17_n_1343) | (mul_34_17_n_2910 & mul_34_17_n_1351));
 assign mul_34_17_n_4554 = ~((mul_34_17_n_1753 & mul_34_17_n_2428) | (mul_34_17_n_2878 & mul_34_17_n_2594));
 assign mul_34_17_n_4553 = ~((mul_34_17_n_1739 & mul_34_17_n_1972) | (mul_34_17_n_2884 & mul_34_17_n_2491));
 assign mul_34_17_n_4552 = ~((mul_34_17_n_669 & mul_34_17_n_1169) | (mul_34_17_n_2916 & mul_34_17_n_1148));
 assign mul_34_17_n_4551 = ~((mul_34_17_n_1745 & mul_34_17_n_2303) | (mul_34_17_n_2888 & mul_34_17_n_2561));
 assign mul_34_17_n_4550 = ((mul_34_17_n_664 | mul_34_17_n_1282) & (mul_34_17_n_11564 | mul_34_17_n_1295));
 assign mul_34_17_n_4549 = ~((mul_34_17_n_679 & mul_34_17_n_911) | (mul_34_17_n_2926 & mul_34_17_n_912));
 assign mul_34_17_n_4548 = ~((mul_34_17_n_1751 & mul_34_17_n_2635) | (mul_34_17_n_2880 & mul_34_17_n_1964));
 assign mul_34_17_n_4547 = ~((mul_34_17_n_665 & mul_34_17_n_1253) | (mul_34_17_n_2912 & mul_34_17_n_1298));
 assign mul_34_17_n_4546 = ~((mul_34_17_n_1753 & mul_34_17_n_1995) | (mul_34_17_n_2878 & mul_34_17_n_2593));
 assign mul_34_17_n_4545 = ~((mul_34_17_n_677 & mul_34_17_n_937) | (mul_34_17_n_2924 & mul_34_17_n_933));
 assign mul_34_17_n_4544 = ~((mul_34_17_n_1735 & mul_34_17_n_2501) | (mul_34_17_n_2896 & mul_34_17_n_2591));
 assign mul_34_17_n_4543 = ~((mul_34_17_n_667 & mul_34_17_n_1202) | (mul_34_17_n_2914 & mul_34_17_n_1214));
 assign mul_34_17_n_4542 = ((mul_34_17_n_1748 | mul_34_17_n_1694) & (mul_34_17_n_11597 | mul_34_17_n_2645));
 assign mul_34_17_n_4541 = ~((mul_34_17_n_688 | mul_34_17_n_902) & (mul_34_17_n_11528 | mul_34_17_n_700));
 assign mul_34_17_n_4540 = ((mul_34_17_n_1750 | mul_34_17_n_2089) & (mul_34_17_n_11612 | mul_34_17_n_2531));
 assign mul_34_17_n_4539 = ((mul_34_17_n_690 | mul_34_17_n_728) & (mul_34_17_n_11525 | mul_34_17_n_702));
 assign mul_34_17_n_4538 = ~((mul_34_17_n_669 & mul_34_17_n_1158) | (mul_34_17_n_2916 & mul_34_17_n_1136));
 assign mul_34_17_n_4537 = ~((mul_34_17_n_1739 & mul_34_17_n_2596) | (mul_34_17_n_2884 & mul_34_17_n_2159));
 assign mul_34_17_n_4536 = ((mul_34_17_n_666 | mul_34_17_n_1185) & (mul_34_17_n_11561 | mul_34_17_n_1238));
 assign mul_34_17_n_4535 = ~((mul_34_17_n_691 & mul_34_17_n_715) | (mul_34_17_n_2936 & mul_34_17_n_729));
 assign mul_34_17_n_4534 = ~((mul_34_17_n_1753 & mul_34_17_n_2590) | (mul_34_17_n_2878 & mul_34_17_n_2359));
 assign mul_34_17_n_4533 = ((mul_34_17_n_655 & mul_34_17_n_1602) | (mul_34_17_n_2902 & mul_34_17_n_1648));
 assign mul_34_17_n_4532 = ~((mul_34_17_n_657 & mul_34_17_n_1584) | (mul_34_17_n_2904 & mul_34_17_n_1523));
 assign mul_34_17_n_4530 = ((mul_34_17_n_1742 | mul_34_17_n_1943) & (mul_34_17_n_11609 | mul_34_17_n_2155));
 assign mul_34_17_n_4529 = ((mul_34_17_n_1756 | mul_34_17_n_1675) & (mul_34_17_n_11582 | mul_34_17_n_1686));
 assign mul_34_17_n_4528 = ((mul_34_17_n_1742 | mul_34_17_n_2592) & (mul_34_17_n_11609 | mul_34_17_n_2371));
 assign mul_34_17_n_4527 = ((mul_34_17_n_672 | mul_34_17_n_1066) & (mul_34_17_n_11552 | mul_34_17_n_1064));
 assign mul_34_17_n_4526 = ~((mul_34_17_n_1743 & mul_34_17_n_2490) | (mul_34_17_n_2882 & mul_34_17_n_2109));
 assign mul_34_17_n_4525 = ((mul_34_17_n_1745 & mul_34_17_n_2382) | (mul_34_17_n_2888 & mul_34_17_n_2502));
 assign mul_34_17_n_4524 = ((mul_34_17_n_1754 | mul_34_17_n_2681) & (mul_34_17_n_11585 | mul_34_17_n_2548));
 assign mul_34_17_n_4523 = ~((mul_34_17_n_675 & mul_34_17_n_976) | (mul_34_17_n_2922 & mul_34_17_n_1001));
 assign mul_34_17_n_4522 = ~((mul_34_17_n_671 & mul_34_17_n_1076) | (mul_34_17_n_2918 & mul_34_17_n_1072));
 assign mul_34_17_n_4520 = ((mul_34_17_n_656 | mul_34_17_n_1551) & (mul_34_17_n_11576 | mul_34_17_n_1568));
 assign mul_34_17_n_4519 = ((mul_34_17_n_1757 & mul_34_17_n_2261) | (mul_34_17_n_2900 & mul_34_17_n_2163));
 assign mul_34_17_n_4518 = ~((mul_34_17_n_673 & mul_34_17_n_1044) | (mul_34_17_n_2920 & mul_34_17_n_1018));
 assign mul_34_17_n_4517 = ~((mul_34_17_n_659 & mul_34_17_n_1459) | (mul_34_17_n_2906 & mul_34_17_n_1504));
 assign mul_34_17_n_4515 = ((mul_34_17_n_1734 | mul_34_17_n_2692) & (mul_34_17_n_11588 | mul_34_17_n_1894));
 assign mul_34_17_n_4513 = ((mul_34_17_n_682 | mul_34_17_n_812) & (mul_34_17_n_11537 | mul_34_17_n_832));
 assign mul_34_17_n_4511 = ((mul_34_17_n_658 | mul_34_17_n_1457) & (mul_34_17_n_11573 | mul_34_17_n_1474));
 assign mul_34_17_n_4509 = ((mul_34_17_n_1748 | mul_34_17_n_2006) & (mul_34_17_n_11597 | mul_34_17_n_2556));
 assign mul_34_17_n_4508 = ~((mul_34_17_n_1741 & mul_34_17_n_2190) | (mul_34_17_n_2886 & mul_34_17_n_2331));
 assign mul_34_17_n_4507 = ~((mul_34_17_n_661 & mul_34_17_n_1433) | (mul_34_17_n_2908 & mul_34_17_n_1384));
 assign mul_34_17_n_4505 = ~((mul_34_17_n_663 & mul_34_17_n_1351) | (mul_34_17_n_2910 & mul_34_17_n_1325));
 assign mul_34_17_n_4504 = ~((mul_34_17_n_1737 & mul_34_17_n_2355) | (mul_34_17_n_2894 & mul_34_17_n_2429));
 assign mul_34_17_n_4503 = ~((mul_34_17_n_1747 & mul_34_17_n_2169) | (mul_34_17_n_11593 & mul_34_17_n_2426));
 assign mul_34_17_n_4501 = ~((mul_34_17_n_1743 & mul_34_17_n_2664) | (mul_34_17_n_2882 & mul_34_17_n_2370));
 assign mul_34_17_n_4500 = ~((mul_34_17_n_1745 & mul_34_17_n_2597) | (mul_34_17_n_2888 & mul_34_17_n_2095));
 assign mul_34_17_n_4499 = ~((mul_34_17_n_687 & mul_34_17_n_743) | (mul_34_17_n_2933 & mul_34_17_n_718));
 assign mul_34_17_n_4498 = ~((mul_34_17_n_1743 & mul_34_17_n_1903) | (mul_34_17_n_2882 & mul_34_17_n_2334));
 assign mul_34_17_n_4496 = ~((mul_34_17_n_671 & mul_34_17_n_1120) | (mul_34_17_n_2918 & mul_34_17_n_1073));
 assign mul_34_17_n_4494 = ~((mul_34_17_n_673 & mul_34_17_n_1051) | (mul_34_17_n_2920 & mul_34_17_n_1016));
 assign mul_34_17_n_4493 = ~((mul_34_17_n_655 & mul_34_17_n_1622) | (mul_34_17_n_2902 & mul_34_17_n_1660));
 assign mul_34_17_n_4492 = ((mul_34_17_n_1755 & mul_34_17_n_2483) | (mul_34_17_n_2898 & mul_34_17_n_2434));
 assign mul_34_17_n_4491 = ~((mul_34_17_n_1753 & mul_34_17_n_2593) | (mul_34_17_n_2878 & mul_34_17_n_2433));
 assign mul_34_17_n_4490 = ~((mul_34_17_n_493 | mul_34_17_n_494) & (mul_34_17_n_2878 | mul_34_17_n_1753));
 assign mul_34_17_n_4488 = ~((mul_34_17_n_1751 & mul_34_17_n_2623) | (mul_34_17_n_2880 & mul_34_17_n_2578));
 assign mul_34_17_n_4487 = ((mul_34_17_n_1757 & mul_34_17_n_2435) | (mul_34_17_n_2900 & mul_34_17_n_1759));
 assign mul_34_17_n_4486 = ((mul_34_17_n_688 | mul_34_17_n_701) & (mul_34_17_n_11528 | mul_34_17_n_936));
 assign mul_34_17_n_4484 = ~((mul_34_17_n_665 & mul_34_17_n_1298) | (mul_34_17_n_2912 & mul_34_17_n_1249));
 assign mul_34_17_n_4483 = ~((mul_34_17_n_673 & mul_34_17_n_1055) | (mul_34_17_n_2920 & mul_34_17_n_1053));
 assign mul_34_17_n_4482 = ~((mul_34_17_n_1749 & mul_34_17_n_1850) | (mul_34_17_n_2890 & mul_34_17_n_2569));
 assign mul_34_17_n_4481 = ~((mul_34_17_n_1757 & mul_34_17_n_1767) | (mul_34_17_n_2900 & mul_34_17_n_1760));
 assign mul_34_17_n_4480 = ~((mul_34_17_n_661 & mul_34_17_n_1437) | (mul_34_17_n_2908 & mul_34_17_n_1441));
 assign mul_34_17_n_4479 = ~((mul_34_17_n_667 & mul_34_17_n_1204) | (mul_34_17_n_2914 & mul_34_17_n_1224));
 assign mul_34_17_n_4478 = ~(mul_34_17_n_3003 | mul_34_17_n_2753);
 assign mul_34_17_n_4477 = ~((mul_34_17_n_667 & mul_34_17_n_1245) | (mul_34_17_n_2914 & mul_34_17_n_1246));
 assign mul_34_17_n_4476 = ~((mul_34_17_n_669 & mul_34_17_n_1148) | (mul_34_17_n_2916 & mul_34_17_n_1147));
 assign mul_34_17_n_4475 = ((mul_34_17_n_1750 | mul_34_17_n_1991) & (mul_34_17_n_11612 | mul_34_17_n_1855));
 assign mul_34_17_n_4474 = ~((mul_34_17_n_1743 & mul_34_17_n_2409) | (mul_34_17_n_2882 & mul_34_17_n_2505));
 assign mul_34_17_n_4473 = ~(mul_34_17_n_3002 | mul_34_17_n_2752);
 assign mul_34_17_n_4472 = ~((mul_34_17_n_661 & mul_34_17_n_1428) | (mul_34_17_n_2908 & mul_34_17_n_1374));
 assign mul_34_17_n_4471 = ~((mul_34_17_n_1743 & mul_34_17_n_1876) | (mul_34_17_n_2882 & mul_34_17_n_2648));
 assign mul_34_17_n_4470 = ~((mul_34_17_n_1757 & mul_34_17_n_1632) | (mul_34_17_n_2900 & mul_34_17_n_828));
 assign mul_34_17_n_4469 = ((mul_34_17_n_676 | mul_34_17_n_924) & (mul_34_17_n_11546 | mul_34_17_n_965));
 assign mul_34_17_n_4468 = ((mul_34_17_n_686 | mul_34_17_n_757) & (mul_34_17_n_11531 | mul_34_17_n_748));
 assign mul_34_17_n_4467 = ~((mul_34_17_n_663 & mul_34_17_n_1344) | (mul_34_17_n_2910 & mul_34_17_n_1334));
 assign mul_34_17_n_4465 = ~((mul_34_17_n_1753 & mul_34_17_n_1840) | (mul_34_17_n_2878 & mul_34_17_n_1993));
 assign mul_34_17_n_4463 = ((mul_34_17_n_1736 | mul_34_17_n_2436) & (mul_34_17_n_11591 | mul_34_17_n_2460));
 assign mul_34_17_n_4462 = ((mul_34_17_n_1748 | mul_34_17_n_2506) & (mul_34_17_n_11597 | mul_34_17_n_2485));
 assign mul_34_17_n_4460 = ~((mul_34_17_n_1741 & mul_34_17_n_2151) | (mul_34_17_n_2886 & mul_34_17_n_1947));
 assign mul_34_17_n_4458 = ~((mul_34_17_n_1757 & mul_34_17_n_2542) | (mul_34_17_n_2900 & mul_34_17_n_1676));
 assign mul_34_17_n_4457 = ((mul_34_17_n_1743 & mul_34_17_n_1956) | (mul_34_17_n_2882 & mul_34_17_n_2468));
 assign mul_34_17_n_4456 = ~(mul_34_17_n_2996 | mul_34_17_n_2751);
 assign mul_34_17_n_4455 = ~((mul_34_17_n_1737 & mul_34_17_n_2611) | (mul_34_17_n_2894 & mul_34_17_n_2278));
 assign mul_34_17_n_4453 = ~((mul_34_17_n_669 & mul_34_17_n_1144) | (mul_34_17_n_2916 & mul_34_17_n_1153));
 assign mul_34_17_n_4452 = ((mul_34_17_n_1736 | mul_34_17_n_2346) & (mul_34_17_n_11591 | mul_34_17_n_2293));
 assign mul_34_17_n_4451 = ~((mul_34_17_n_655 & mul_34_17_n_1662) | (mul_34_17_n_2902 & mul_34_17_n_1595));
 assign mul_34_17_n_4450 = ((mul_34_17_n_654 | mul_34_17_n_1590) & (mul_34_17_n_11579 | mul_34_17_n_1640));
 assign mul_34_17_n_4449 = ~((mul_34_17_n_1747 & mul_34_17_n_2276) | (mul_34_17_n_11593 & mul_34_17_n_2570));
 assign mul_34_17_n_4448 = ~((mul_34_17_n_673 & mul_34_17_n_1046) | (mul_34_17_n_2920 & mul_34_17_n_1033));
 assign mul_34_17_n_4446 = ((mul_34_17_n_654 | mul_34_17_n_1599) & (mul_34_17_n_11579 | mul_34_17_n_1636));
 assign mul_34_17_n_4445 = ~((mul_34_17_n_663 & mul_34_17_n_1357) | (mul_34_17_n_2910 & mul_34_17_n_1371));
 assign mul_34_17_n_4444 = ~((mul_34_17_n_1739 & mul_34_17_n_2309) | (mul_34_17_n_2884 & mul_34_17_n_2666));
 assign mul_34_17_n_4443 = ~((mul_34_17_n_655 & mul_34_17_n_1646) | (mul_34_17_n_2902 & mul_34_17_n_1664));
 assign mul_34_17_n_4442 = ((mul_34_17_n_671 & mul_34_17_n_1106) | (mul_34_17_n_2918 & mul_34_17_n_1083));
 assign mul_34_17_n_4441 = ((mul_34_17_n_688 | mul_34_17_n_703) & (mul_34_17_n_11528 | mul_34_17_n_726));
 assign mul_34_17_n_4439 = ((mul_34_17_n_688 | mul_34_17_n_936) & (mul_34_17_n_11528 | mul_34_17_n_692));
 assign mul_34_17_n_4437 = ~((mul_34_17_n_665 & mul_34_17_n_1283) | (mul_34_17_n_2912 & mul_34_17_n_1297));
 assign mul_34_17_n_4436 = ~((mul_34_17_n_657 & mul_34_17_n_1559) | (mul_34_17_n_2904 & mul_34_17_n_1567));
 assign mul_34_17_n_4434 = ~((mul_34_17_n_681 & mul_34_17_n_871) | (mul_34_17_n_2928 & mul_34_17_n_838));
 assign mul_34_17_n_4432 = ~((mul_34_17_n_691 & mul_34_17_n_705) | (mul_34_17_n_2936 & mul_34_17_n_742));
 assign mul_34_17_n_4430 = ~((mul_34_17_n_661 & mul_34_17_n_1384) | (mul_34_17_n_2908 & mul_34_17_n_1426));
 assign mul_34_17_n_4429 = ((mul_34_17_n_684 | mul_34_17_n_782) & (mul_34_17_n_11534 | mul_34_17_n_784));
 assign mul_34_17_n_4427 = ~((mul_34_17_n_685 & mul_34_17_n_789) | (mul_34_17_n_2931 & mul_34_17_n_794));
 assign mul_34_17_n_4426 = ~((mul_34_17_n_661 & mul_34_17_n_1394) | (mul_34_17_n_2908 & mul_34_17_n_1408));
 assign mul_34_17_n_4424 = ~((mul_34_17_n_677 & mul_34_17_n_939) | (mul_34_17_n_2924 & mul_34_17_n_960));
 assign mul_34_17_n_4423 = ~((mul_34_17_n_665 & mul_34_17_n_1277) | (mul_34_17_n_2912 & mul_34_17_n_1289));
 assign mul_34_17_n_4422 = ((mul_34_17_n_671 & mul_34_17_n_1079) | (mul_34_17_n_2918 & mul_34_17_n_1099));
 assign mul_34_17_n_4420 = ((mul_34_17_n_682 | mul_34_17_n_832) & (mul_34_17_n_11537 | mul_34_17_n_824));
 assign mul_34_17_n_4418 = ~((mul_34_17_n_669 & mul_34_17_n_1147) | (mul_34_17_n_2916 & mul_34_17_n_1132));
 assign mul_34_17_n_4417 = ~((mul_34_17_n_671 & mul_34_17_n_1096) | (mul_34_17_n_2918 & mul_34_17_n_1120));
 assign mul_34_17_n_4416 = ~((mul_34_17_n_685 & mul_34_17_n_788) | (mul_34_17_n_2931 & mul_34_17_n_777));
 assign mul_34_17_n_4415 = ((mul_34_17_n_682 | mul_34_17_n_830) & (mul_34_17_n_11537 | mul_34_17_n_833));
 assign mul_34_17_n_4414 = ((mul_34_17_n_682 | mul_34_17_n_815) & (mul_34_17_n_11537 | mul_34_17_n_812));
 assign mul_34_17_n_4413 = ((mul_34_17_n_664 | mul_34_17_n_1305) & (mul_34_17_n_11564 | mul_34_17_n_1307));
 assign mul_34_17_n_4412 = ~(mul_34_17_n_2864 ^ mul_34_17_n_2969);
 assign mul_34_17_n_4411 = ~((mul_34_17_n_665 & mul_34_17_n_1290) | (mul_34_17_n_2912 & mul_34_17_n_1277));
 assign mul_34_17_n_4410 = ~((mul_34_17_n_661 & mul_34_17_n_1438) | (mul_34_17_n_2908 & mul_34_17_n_1418));
 assign mul_34_17_n_4409 = ~((mul_34_17_n_1743 & mul_34_17_n_1689) | (mul_34_17_n_2882 & mul_34_17_n_2497));
 assign mul_34_17_n_4408 = ((mul_34_17_n_1734 | mul_34_17_n_1892) & (mul_34_17_n_11588 | mul_34_17_n_2688));
 assign mul_34_17_n_4407 = ~((mul_34_17_n_685 & mul_34_17_n_795) | (mul_34_17_n_2931 & mul_34_17_n_783));
 assign mul_34_17_n_4406 = ~((mul_34_17_n_661 & mul_34_17_n_1409) | (mul_34_17_n_2908 & mul_34_17_n_1435));
 assign mul_34_17_n_4405 = ~((mul_34_17_n_663 & mul_34_17_n_1311) | (mul_34_17_n_2910 & mul_34_17_n_1369));
 assign mul_34_17_n_4404 = ~((mul_34_17_n_1753 & mul_34_17_n_2433) | (mul_34_17_n_2878 & mul_34_17_n_2287));
 assign mul_34_17_n_4403 = ~((mul_34_17_n_682 | mul_34_17_n_803) & (mul_34_17_n_11537 | mul_34_17_n_822));
 assign mul_34_17_n_4402 = ~((mul_34_17_n_671 & mul_34_17_n_1087) | (mul_34_17_n_2918 & mul_34_17_n_1086));
 assign mul_34_17_n_4401 = ~((mul_34_17_n_671 & mul_34_17_n_1073) | (mul_34_17_n_2918 & mul_34_17_n_1125));
 assign mul_34_17_n_4400 = ((mul_34_17_n_680 | mul_34_17_n_850) & (mul_34_17_n_11540 | mul_34_17_n_836));
 assign mul_34_17_n_4399 = ~((mul_34_17_n_1737 & mul_34_17_n_1897) | (mul_34_17_n_2894 & mul_34_17_n_2546));
 assign mul_34_17_n_4398 = ~((mul_34_17_n_1749 & mul_34_17_n_2532) | (mul_34_17_n_2890 & mul_34_17_n_2415));
 assign mul_34_17_n_4397 = ((mul_34_17_n_1753 & mul_34_17_n_1993) | (mul_34_17_n_2878 & mul_34_17_n_2397));
 assign mul_34_17_n_4396 = ((mul_34_17_n_680 | mul_34_17_n_859) & (mul_34_17_n_11540 | mul_34_17_n_844));
 assign mul_34_17_n_4395 = ~((mul_34_17_n_669 & mul_34_17_n_1153) | (mul_34_17_n_2916 & mul_34_17_n_1151));
 assign mul_34_17_n_4394 = ~((mul_34_17_n_657 & mul_34_17_n_1586) | (mul_34_17_n_2904 & mul_34_17_n_1533));
 assign mul_34_17_n_4393 = ~((mul_34_17_n_687 & mul_34_17_n_1589) | (mul_34_17_n_2933 & mul_34_17_n_758));
 assign mul_34_17_n_4392 = ~((mul_34_17_n_659 & mul_34_17_n_1448) | (mul_34_17_n_2906 & mul_34_17_n_1509));
 assign mul_34_17_n_4391 = ~(mul_34_17_n_2941 ^ mul_34_17_n_2863);
 assign mul_34_17_n_4389 = ~((mul_34_17_n_1745 & mul_34_17_n_2124) | (mul_34_17_n_2888 & mul_34_17_n_2482));
 assign mul_34_17_n_4388 = ~((mul_34_17_n_657 & mul_34_17_n_1577) | (mul_34_17_n_2904 & mul_34_17_n_1585));
 assign mul_34_17_n_4387 = ~((mul_34_17_n_669 & mul_34_17_n_1141) | (mul_34_17_n_2916 & mul_34_17_n_1179));
 assign mul_34_17_n_4386 = ((mul_34_17_n_1752 | mul_34_17_n_2410) & (mul_34_17_n_11615 | mul_34_17_n_2650));
 assign mul_34_17_n_4385 = ~((mul_34_17_n_655 & mul_34_17_n_1619) | (mul_34_17_n_2902 & mul_34_17_n_1613));
 assign mul_34_17_n_4383 = ~((mul_34_17_n_677 & mul_34_17_n_925) | (mul_34_17_n_2924 & mul_34_17_n_946));
 assign mul_34_17_n_4382 = ((mul_34_17_n_676 | mul_34_17_n_962) & (mul_34_17_n_11546 | mul_34_17_n_924));
 assign mul_34_17_n_4380 = ~((mul_34_17_n_675 & mul_34_17_n_1011) | (mul_34_17_n_2922 & mul_34_17_n_981));
 assign mul_34_17_n_4379 = ((mul_34_17_n_674 | mul_34_17_n_1004) & (mul_34_17_n_11549 | mul_34_17_n_1013));
 assign mul_34_17_n_4378 = ((mul_34_17_n_1746 | mul_34_17_n_2367) & (mul_34_17_n_11648 | mul_34_17_n_2585));
 assign mul_34_17_n_4377 = ~((mul_34_17_n_1751 & mul_34_17_n_2626) | (mul_34_17_n_2880 & mul_34_17_n_2200));
 assign mul_34_17_n_4376 = ~((mul_34_17_n_1757 & mul_34_17_n_1685) | (mul_34_17_n_2900 & mul_34_17_n_2097));
 assign mul_34_17_n_4375 = ~((mul_34_17_n_1751 & mul_34_17_n_2644) | (mul_34_17_n_2880 & mul_34_17_n_2134));
 assign mul_34_17_n_4374 = ~((mul_34_17_n_659 & mul_34_17_n_1460) | (mul_34_17_n_2906 & mul_34_17_n_1477));
 assign mul_34_17_n_4373 = ~((mul_34_17_n_665 & mul_34_17_n_1272) | (mul_34_17_n_2912 & mul_34_17_n_1257));
 assign mul_34_17_n_4372 = ~(mul_34_17_n_2870 ^ mul_34_17_n_2952);
 assign mul_34_17_n_4371 = ~((mul_34_17_n_1743 & mul_34_17_n_2612) | (mul_34_17_n_2882 & mul_34_17_n_1966));
 assign mul_34_17_n_4369 = ~((mul_34_17_n_665 & mul_34_17_n_1257) | (mul_34_17_n_2912 & mul_34_17_n_1306));
 assign mul_34_17_n_4368 = ((mul_34_17_n_655 & mul_34_17_n_1605) | (mul_34_17_n_2902 & mul_34_17_n_1606));
 assign mul_34_17_n_4366 = ((mul_34_17_n_688 | mul_34_17_n_709) & (mul_34_17_n_11528 | mul_34_17_n_1266));
 assign mul_34_17_n_4365 = ~((mul_34_17_n_1739 & mul_34_17_n_2373) | (mul_34_17_n_2884 & mul_34_17_n_1972));
 assign mul_34_17_n_4364 = ~((mul_34_17_n_663 & mul_34_17_n_1324) | (mul_34_17_n_2910 & mul_34_17_n_1329));
 assign mul_34_17_n_4363 = ~((mul_34_17_n_661 & mul_34_17_n_1377) | (mul_34_17_n_2908 & mul_34_17_n_1434));
 assign mul_34_17_n_4362 = ~((mul_34_17_n_1751 & mul_34_17_n_1960) | (mul_34_17_n_2880 & mul_34_17_n_2623));
 assign mul_34_17_n_4361 = ((mul_34_17_n_676 | mul_34_17_n_950) & (mul_34_17_n_11546 | mul_34_17_n_931));
 assign mul_34_17_n_4360 = ((mul_34_17_n_1756 | mul_34_17_n_1958) & (mul_34_17_n_11582 | mul_34_17_n_1279));
 assign mul_34_17_n_4359 = ((mul_34_17_n_664 | mul_34_17_n_1302) & (mul_34_17_n_11564 | mul_34_17_n_1274));
 assign mul_34_17_n_4358 = ~((mul_34_17_n_671 & mul_34_17_n_1108) | (mul_34_17_n_2918 & mul_34_17_n_1102));
 assign mul_34_17_n_4357 = ((mul_34_17_n_1734 | mul_34_17_n_2683) & (mul_34_17_n_11588 | mul_34_17_n_2186));
 assign mul_34_17_n_4356 = ~((mul_34_17_n_681 & mul_34_17_n_856) | (mul_34_17_n_2928 & mul_34_17_n_860));
 assign mul_34_17_n_4355 = ~((mul_34_17_n_657 & mul_34_17_n_1555) | (mul_34_17_n_2904 & mul_34_17_n_1560));
 assign mul_34_17_n_4354 = ~((mul_34_17_n_687 & mul_34_17_n_1385) | (mul_34_17_n_2933 & mul_34_17_n_1589));
 assign mul_34_17_n_4353 = ~((mul_34_17_n_1753 & mul_34_17_n_2114) | (mul_34_17_n_2878 & mul_34_17_n_2498));
 assign mul_34_17_n_4352 = ~((mul_34_17_n_1741 & mul_34_17_n_2193) | (mul_34_17_n_2886 & mul_34_17_n_2621));
 assign mul_34_17_n_4351 = ((mul_34_17_n_1748 | mul_34_17_n_2271) & (mul_34_17_n_11597 | mul_34_17_n_2671));
 assign mul_34_17_n_4349 = ~((mul_34_17_n_1747 & mul_34_17_n_2467) | (mul_34_17_n_11593 & mul_34_17_n_2174));
 assign mul_34_17_n_4348 = ~((mul_34_17_n_657 & mul_34_17_n_1560) | (mul_34_17_n_2904 & mul_34_17_n_1573));
 assign mul_34_17_n_4347 = ((mul_34_17_n_688 | mul_34_17_n_842) & (mul_34_17_n_11528 | mul_34_17_n_769));
 assign mul_34_17_n_4346 = ((mul_34_17_n_656 | mul_34_17_n_1553) & (mul_34_17_n_11576 | mul_34_17_n_1549));
 assign mul_34_17_n_4345 = ~((mul_34_17_n_667 & mul_34_17_n_1212) | (mul_34_17_n_2914 & mul_34_17_n_1195));
 assign mul_34_17_n_4344 = ((mul_34_17_n_1734 | mul_34_17_n_2264) & (mul_34_17_n_11588 | mul_34_17_n_2441));
 assign mul_34_17_n_4342 = ~((mul_34_17_n_1757 & mul_34_17_n_2163) | (mul_34_17_n_2900 & mul_34_17_n_1003));
 assign mul_34_17_n_4341 = ~((mul_34_17_n_663 & mul_34_17_n_1367) | (mul_34_17_n_2910 & mul_34_17_n_1343));
 assign mul_34_17_n_4340 = ((mul_34_17_n_666 | mul_34_17_n_1220) & (mul_34_17_n_11561 | mul_34_17_n_1222));
 assign mul_34_17_n_4338 = ~((mul_34_17_n_1751 & mul_34_17_n_2043) | (mul_34_17_n_2880 & mul_34_17_n_2086));
 assign mul_34_17_n_4336 = ~((mul_34_17_n_665 & mul_34_17_n_1249) | (mul_34_17_n_2912 & mul_34_17_n_1261));
 assign mul_34_17_n_4335 = ~((mul_34_17_n_1743 & mul_34_17_n_1863) | (mul_34_17_n_2882 & mul_34_17_n_2424));
 assign mul_34_17_n_4334 = ~(mul_34_17_n_2997 | mul_34_17_n_2747);
 assign mul_34_17_n_4332 = ~((mul_34_17_n_1747 & mul_34_17_n_2381) | (mul_34_17_n_11593 & mul_34_17_n_2691));
 assign mul_34_17_n_4331 = ((mul_34_17_n_1748 | mul_34_17_n_2509) & (mul_34_17_n_11597 | mul_34_17_n_2237));
 assign mul_34_17_n_4329 = ~((mul_34_17_n_1755 & mul_34_17_n_2434) | (mul_34_17_n_2898 & mul_34_17_n_2447));
 assign mul_34_17_n_4328 = ((mul_34_17_n_654 | mul_34_17_n_1627) & (mul_34_17_n_11579 | mul_34_17_n_1645));
 assign mul_34_17_n_4326 = ~((mul_34_17_n_1747 & mul_34_17_n_1886) | (mul_34_17_n_11593 & mul_34_17_n_1870));
 assign mul_34_17_n_4325 = ((mul_34_17_n_659 & mul_34_17_n_1472) | (mul_34_17_n_2906 & mul_34_17_n_1516));
 assign mul_34_17_n_4324 = ~((mul_34_17_n_657 & mul_34_17_n_1541) | (mul_34_17_n_2904 & mul_34_17_n_1577));
 assign mul_34_17_n_4323 = ((mul_34_17_n_661 & mul_34_17_n_1396) | (mul_34_17_n_2908 & mul_34_17_n_1400));
 assign mul_34_17_n_4321 = ~((mul_34_17_n_1735 & mul_34_17_n_2379) | (mul_34_17_n_2896 & mul_34_17_n_2528));
 assign mul_34_17_n_4320 = ((mul_34_17_n_657 & mul_34_17_n_1535) | (mul_34_17_n_2904 & mul_34_17_n_1554));
 assign mul_34_17_n_4318 = ~((mul_34_17_n_1739 & mul_34_17_n_1957) | (mul_34_17_n_2884 & mul_34_17_n_1860));
 assign mul_34_17_n_4317 = ((mul_34_17_n_1751 & mul_34_17_n_2047) | (mul_34_17_n_2880 & mul_34_17_n_2527));
 assign mul_34_17_n_4316 = ((mul_34_17_n_1753 & mul_34_17_n_1873) | (mul_34_17_n_2878 & mul_34_17_n_2540));
 assign mul_34_17_n_4315 = ((mul_34_17_n_682 | mul_34_17_n_821) & (mul_34_17_n_11537 | mul_34_17_n_804));
 assign mul_34_17_n_4314 = ~(mul_34_17_n_2998 | mul_34_17_n_2754);
 assign mul_34_17_n_4313 = ~((mul_34_17_n_1743 & mul_34_17_n_2488) | (mul_34_17_n_2882 & mul_34_17_n_1871));
 assign mul_34_17_n_4312 = ~((mul_34_17_n_675 & mul_34_17_n_981) | (mul_34_17_n_2922 & mul_34_17_n_1012));
 assign mul_34_17_n_4310 = ~((mul_34_17_n_1745 & mul_34_17_n_2651) | (mul_34_17_n_2888 & mul_34_17_n_2273));
 assign mul_34_17_n_4309 = ~((mul_34_17_n_679 & mul_34_17_n_892) | (mul_34_17_n_2926 & mul_34_17_n_910));
 assign mul_34_17_n_4308 = ((mul_34_17_n_685 & mul_34_17_n_785) | (mul_34_17_n_2931 & mul_34_17_n_796));
 assign mul_34_17_n_4307 = ~((mul_34_17_n_1749 & mul_34_17_n_2247) | (mul_34_17_n_2890 & mul_34_17_n_1848));
 assign mul_34_17_n_4305 = ((mul_34_17_n_1740 | mul_34_17_n_2038) & (mul_34_17_n_11603 | mul_34_17_n_1933));
 assign mul_34_17_n_4303 = ((mul_34_17_n_666 | mul_34_17_n_1225) & (mul_34_17_n_11561 | mul_34_17_n_1220));
 assign mul_34_17_n_4302 = ((mul_34_17_n_665 & mul_34_17_n_1251) | (mul_34_17_n_2912 & mul_34_17_n_1258));
 assign mul_34_17_n_4300 = ~((mul_34_17_n_673 & mul_34_17_n_1065) | (mul_34_17_n_2920 & mul_34_17_n_1061));
 assign mul_34_17_n_4299 = ~((mul_34_17_n_1737 & mul_34_17_n_1866) | (mul_34_17_n_2894 & mul_34_17_n_2427));
 assign mul_34_17_n_4298 = ((mul_34_17_n_664 | mul_34_17_n_1262) & (mul_34_17_n_11564 | mul_34_17_n_1302));
 assign mul_34_17_n_4297 = ((mul_34_17_n_1742 | mul_34_17_n_1988) & (mul_34_17_n_11609 | mul_34_17_n_2298));
 assign mul_34_17_n_4296 = ((mul_34_17_n_662 | mul_34_17_n_1316) & (mul_34_17_n_11567 | mul_34_17_n_1323));
 assign mul_34_17_n_4295 = ~((mul_34_17_n_1745 & mul_34_17_n_2587) | (mul_34_17_n_2888 & mul_34_17_n_2119));
 assign mul_34_17_n_4293 = ~((mul_34_17_n_1739 & mul_34_17_n_2639) | (mul_34_17_n_2884 & mul_34_17_n_2113));
 assign mul_34_17_n_4292 = ~((mul_34_17_n_1735 & mul_34_17_n_2082) | (mul_34_17_n_2896 & mul_34_17_n_2690));
 assign mul_34_17_n_4291 = ~((mul_34_17_n_1741 & mul_34_17_n_2418) | (mul_34_17_n_2886 & mul_34_17_n_2378));
 assign mul_34_17_n_4290 = ((mul_34_17_n_659 & mul_34_17_n_1490) | (mul_34_17_n_2906 & mul_34_17_n_1453));
 assign mul_34_17_n_4289 = ~((mul_34_17_n_1755 & mul_34_17_n_1843) | (mul_34_17_n_2898 & mul_34_17_n_2059));
 assign mul_34_17_n_4288 = ~((mul_34_17_n_1749 & mul_34_17_n_2210) | (mul_34_17_n_2890 & mul_34_17_n_1862));
 assign mul_34_17_n_4286 = ~((mul_34_17_n_1751 & mul_34_17_n_2063) | (mul_34_17_n_2880 & mul_34_17_n_2225));
 assign mul_34_17_n_4285 = ~((mul_34_17_n_673 & mul_34_17_n_1014) | (mul_34_17_n_2920 & mul_34_17_n_1049));
 assign mul_34_17_n_4284 = ((mul_34_17_n_1739 & mul_34_17_n_2130) | (mul_34_17_n_2884 & mul_34_17_n_2389));
 assign mul_34_17_n_4283 = ~((mul_34_17_n_1735 & mul_34_17_n_2308) | (mul_34_17_n_2896 & mul_34_17_n_2513));
 assign mul_34_17_n_4282 = ~(mul_34_17_n_2874 ^ mul_34_17_n_2950);
 assign mul_34_17_n_4281 = ~((mul_34_17_n_663 & mul_34_17_n_1346) | (mul_34_17_n_2910 & mul_34_17_n_1359));
 assign mul_34_17_n_4280 = ~((mul_34_17_n_1735 & mul_34_17_n_2565) | (mul_34_17_n_2896 & mul_34_17_n_2501));
 assign mul_34_17_n_4279 = ~((mul_34_17_n_1737 & mul_34_17_n_2573) | (mul_34_17_n_2894 & mul_34_17_n_2056));
 assign mul_34_17_n_4278 = ~((mul_34_17_n_1745 & mul_34_17_n_2318) | (mul_34_17_n_2888 & mul_34_17_n_2018));
 assign mul_34_17_n_4277 = ((mul_34_17_n_661 & mul_34_17_n_1442) | (mul_34_17_n_2908 & mul_34_17_n_1413));
 assign mul_34_17_n_4275 = ~((mul_34_17_n_1749 & mul_34_17_n_1994) | (mul_34_17_n_2890 & mul_34_17_n_2375));
 assign mul_34_17_n_4274 = ~((mul_34_17_n_1743 & mul_34_17_n_2648) | (mul_34_17_n_2882 & mul_34_17_n_1903));
 assign mul_34_17_n_4273 = ~((mul_34_17_n_657 & mul_34_17_n_1583) | (mul_34_17_n_2904 & mul_34_17_n_1578));
 assign mul_34_17_n_4272 = ~((mul_34_17_n_669 & mul_34_17_n_1165) | (mul_34_17_n_2916 & mul_34_17_n_1160));
 assign mul_34_17_n_4270 = ((mul_34_17_n_688 | mul_34_17_n_1200) & (mul_34_17_n_11528 | mul_34_17_n_694));
 assign mul_34_17_n_4269 = ((mul_34_17_n_682 | mul_34_17_n_806) & (mul_34_17_n_11537 | mul_34_17_n_817));
 assign mul_34_17_n_4268 = ~((mul_34_17_n_1749 & mul_34_17_n_2486) | (mul_34_17_n_2890 & mul_34_17_n_2295));
 assign mul_34_17_n_4266 = ~((mul_34_17_n_1751 & mul_34_17_n_2200) | (mul_34_17_n_2880 & mul_34_17_n_2213));
 assign mul_34_17_n_4264 = ~((mul_34_17_n_1745 & mul_34_17_n_2686) | (mul_34_17_n_2888 & mul_34_17_n_2124));
 assign mul_34_17_n_4263 = ~((mul_34_17_n_1751 & mul_34_17_n_2350) | (mul_34_17_n_2880 & mul_34_17_n_2312));
 assign mul_34_17_n_4262 = ~((mul_34_17_n_671 & mul_34_17_n_1085) | (mul_34_17_n_2918 & mul_34_17_n_1122));
 assign mul_34_17_n_4260 = ~((mul_34_17_n_1745 & mul_34_17_n_2636) | (mul_34_17_n_2888 & mul_34_17_n_2035));
 assign mul_34_17_n_4259 = ((mul_34_17_n_1741 & mul_34_17_n_2568) | (mul_34_17_n_2886 & mul_34_17_n_2476));
 assign mul_34_17_n_4258 = ~((mul_34_17_n_1755 & mul_34_17_n_2446) | (mul_34_17_n_2898 & mul_34_17_n_1951));
 assign mul_34_17_n_4257 = ~((mul_34_17_n_1741 & mul_34_17_n_2632) | (mul_34_17_n_2886 & mul_34_17_n_2141));
 assign mul_34_17_n_4255 = ((mul_34_17_n_1753 & mul_34_17_n_2338) | (mul_34_17_n_2878 & mul_34_17_n_1877));
 assign mul_34_17_n_4254 = ((mul_34_17_n_1745 & mul_34_17_n_2228) | (mul_34_17_n_2888 & mul_34_17_n_2518));
 assign mul_34_17_n_4253 = ~((mul_34_17_n_1737 & mul_34_17_n_2631) | (mul_34_17_n_2894 & mul_34_17_n_2244));
 assign mul_34_17_n_4252 = ~((mul_34_17_n_663 & mul_34_17_n_1362) | (mul_34_17_n_2910 & mul_34_17_n_1308));
 assign mul_34_17_n_4251 = ~((mul_34_17_n_1753 & mul_34_17_n_2260) | (mul_34_17_n_2878 & mul_34_17_n_2680));
 assign mul_34_17_n_4250 = ((mul_34_17_n_1747 & mul_34_17_n_2423) | (mul_34_17_n_11593 & mul_34_17_n_2007));
 assign mul_34_17_n_4249 = ((mul_34_17_n_1741 & mul_34_17_n_2378) | (mul_34_17_n_2886 & mul_34_17_n_2451));
 assign mul_34_17_n_4248 = ~(mul_34_17_n_2873 ^ mul_34_17_n_2967);
 assign mul_34_17_n_4247 = ((mul_34_17_n_671 & mul_34_17_n_1099) | (mul_34_17_n_2918 & mul_34_17_n_1118));
 assign mul_34_17_n_4245 = ((mul_34_17_n_1738 | mul_34_17_n_2112) & (mul_34_17_n_11606 | mul_34_17_n_2563));
 assign mul_34_17_n_4244 = ~(mul_34_17_n_3000 | mul_34_17_n_2750);
 assign mul_34_17_n_4242 = ~((mul_34_17_n_1735 & mul_34_17_n_2694) | (mul_34_17_n_2896 & mul_34_17_n_2630));
 assign mul_34_17_n_4241 = ((mul_34_17_n_1739 & mul_34_17_n_2491) | (mul_34_17_n_2884 & mul_34_17_n_1971));
 assign mul_34_17_n_4239 = ~((mul_34_17_n_1757 & mul_34_17_n_1111) | (mul_34_17_n_2900 & mul_34_17_n_1063));
 assign mul_34_17_n_4238 = ((mul_34_17_n_665 & mul_34_17_n_1261) | (mul_34_17_n_2912 & mul_34_17_n_1287));
 assign mul_34_17_n_4237 = ((mul_34_17_n_667 & mul_34_17_n_1242) | (mul_34_17_n_2914 & mul_34_17_n_1240));
 assign mul_34_17_n_4236 = ~((mul_34_17_n_685 & mul_34_17_n_776) | (mul_34_17_n_2931 & mul_34_17_n_781));
 assign mul_34_17_n_4235 = ~((mul_34_17_n_659 & mul_34_17_n_1495) | (mul_34_17_n_2906 & mul_34_17_n_1455));
 assign mul_34_17_n_4234 = ((mul_34_17_n_1742 | mul_34_17_n_1965) & (mul_34_17_n_11609 | mul_34_17_n_2304));
 assign mul_34_17_n_4233 = ~((mul_34_17_n_1741 & mul_34_17_n_2673) | (mul_34_17_n_2886 & mul_34_17_n_1953));
 assign mul_34_17_n_4231 = ~((mul_34_17_n_663 & mul_34_17_n_1336) | (mul_34_17_n_2910 & mul_34_17_n_1362));
 assign mul_34_17_n_4230 = ~((mul_34_17_n_1739 & mul_34_17_n_1934) | (mul_34_17_n_2884 & mul_34_17_n_2687));
 assign mul_34_17_n_4229 = ((mul_34_17_n_663 & mul_34_17_n_1369) | (mul_34_17_n_2910 & mul_34_17_n_1367));
 assign mul_34_17_n_4228 = ~((mul_34_17_n_675 & mul_34_17_n_990) | (mul_34_17_n_2922 & mul_34_17_n_996));
 assign mul_34_17_n_4227 = ((mul_34_17_n_1743 & mul_34_17_n_2345) | (mul_34_17_n_2882 & mul_34_17_n_2454));
 assign mul_34_17_n_4226 = ((mul_34_17_n_670 | mul_34_17_n_1069) & (mul_34_17_n_11555 | mul_34_17_n_1092));
 assign mul_34_17_n_4225 = ((mul_34_17_n_663 & mul_34_17_n_1354) | (mul_34_17_n_2910 & mul_34_17_n_1332));
 assign mul_34_17_n_4224 = ~((mul_34_17_n_1749 & mul_34_17_n_2432) | (mul_34_17_n_2890 & mul_34_17_n_2268));
 assign mul_34_17_n_4223 = ~((mul_34_17_n_665 & mul_34_17_n_1286) | (mul_34_17_n_2912 & mul_34_17_n_1268));
 assign mul_34_17_n_4222 = ((mul_34_17_n_681 & mul_34_17_n_861) | (mul_34_17_n_2928 & mul_34_17_n_835));
 assign mul_34_17_n_4221 = ((mul_34_17_n_658 | mul_34_17_n_1503) & (mul_34_17_n_11573 | mul_34_17_n_1489));
 assign mul_34_17_n_4220 = ~(mul_34_17_n_2876 ^ mul_34_17_n_2964);
 assign mul_34_17_n_4219 = ((mul_34_17_n_659 & mul_34_17_n_1487) | (mul_34_17_n_2906 & mul_34_17_n_1497));
 assign mul_34_17_n_4218 = ((mul_34_17_n_1754 | mul_34_17_n_2154) & (mul_34_17_n_11585 | mul_34_17_n_2026));
 assign mul_34_17_n_4217 = ~((mul_34_17_n_1745 & mul_34_17_n_2463) | (mul_34_17_n_2888 & mul_34_17_n_2138));
 assign mul_34_17_n_4216 = ~((mul_34_17_n_1755 & mul_34_17_n_2088) | (mul_34_17_n_2898 & mul_34_17_n_2662));
 assign mul_34_17_n_4215 = ~((mul_34_17_n_661 & mul_34_17_n_1406) | (mul_34_17_n_2908 & mul_34_17_n_1445));
 assign mul_34_17_n_4214 = ~((mul_34_17_n_679 & mul_34_17_n_888) | (mul_34_17_n_2926 & mul_34_17_n_909));
 assign mul_34_17_n_4213 = ((mul_34_17_n_667 & mul_34_17_n_1197) | (mul_34_17_n_2914 & mul_34_17_n_1186));
 assign mul_34_17_n_4212 = ~((mul_34_17_n_1755 & mul_34_17_n_2662) | (mul_34_17_n_2898 & mul_34_17_n_2668));
 assign mul_34_17_n_4211 = ~((mul_34_17_n_691 & mul_34_17_n_754) | (mul_34_17_n_2936 & mul_34_17_n_732));
 assign mul_34_17_n_4210 = ((mul_34_17_n_677 & mul_34_17_n_945) | (mul_34_17_n_2924 & mul_34_17_n_940));
 assign mul_34_17_n_4209 = ~((mul_34_17_n_655 & mul_34_17_n_1661) | (mul_34_17_n_2902 & mul_34_17_n_1662));
 assign mul_34_17_n_4208 = ((mul_34_17_n_675 & mul_34_17_n_1012) | (mul_34_17_n_2922 & mul_34_17_n_977));
 assign mul_34_17_n_4207 = ~((mul_34_17_n_1747 & mul_34_17_n_2617) | (mul_34_17_n_11593 & mul_34_17_n_2281));
 assign mul_34_17_n_4206 = ~((mul_34_17_n_1749 & mul_34_17_n_2575) | (mul_34_17_n_2890 & mul_34_17_n_2576));
 assign mul_34_17_n_4205 = ~((mul_34_17_n_1753 & mul_34_17_n_2620) | (mul_34_17_n_2878 & mul_34_17_n_1978));
 assign mul_34_17_n_4204 = ~((mul_34_17_n_673 & mul_34_17_n_1018) | (mul_34_17_n_2920 & mul_34_17_n_1043));
 assign mul_34_17_n_4202 = ((mul_34_17_n_654 | mul_34_17_n_1643) & (mul_34_17_n_11579 | mul_34_17_n_1647));
 assign mul_34_17_n_4201 = ~((mul_34_17_n_1741 & mul_34_17_n_2473) | (mul_34_17_n_2886 & mul_34_17_n_2515));
 assign mul_34_17_n_4199 = ~((mul_34_17_n_1755 & mul_34_17_n_2649) | (mul_34_17_n_2898 & mul_34_17_n_2670));
 assign mul_34_17_n_4198 = ((mul_34_17_n_1739 & mul_34_17_n_1860) | (mul_34_17_n_2884 & mul_34_17_n_2586));
 assign mul_34_17_n_4197 = ((mul_34_17_n_1749 & mul_34_17_n_1848) | (mul_34_17_n_2890 & mul_34_17_n_1890));
 assign mul_34_17_n_4196 = ~((mul_34_17_n_1739 & mul_34_17_n_2106) | (mul_34_17_n_2884 & mul_34_17_n_2543));
 assign mul_34_17_n_4195 = ~((mul_34_17_n_1741 & mul_34_17_n_2621) | (mul_34_17_n_2886 & mul_34_17_n_2190));
 assign mul_34_17_n_4194 = ((mul_34_17_n_674 | mul_34_17_n_985) & (mul_34_17_n_11549 | mul_34_17_n_992));
 assign mul_34_17_n_4193 = ~((mul_34_17_n_661 & mul_34_17_n_1391) | (mul_34_17_n_2908 & mul_34_17_n_1410));
 assign mul_34_17_n_4191 = ~((mul_34_17_n_677 & mul_34_17_n_946) | (mul_34_17_n_2924 & mul_34_17_n_945));
 assign mul_34_17_n_4190 = ~((mul_34_17_n_1735 & mul_34_17_n_2659) | (mul_34_17_n_2896 & mul_34_17_n_2070));
 assign mul_34_17_n_4189 = ~((mul_34_17_n_1737 & mul_34_17_n_1977) | (mul_34_17_n_2894 & mul_34_17_n_2611));
 assign mul_34_17_n_4187 = ~((mul_34_17_n_670 | mul_34_17_n_1090) & (mul_34_17_n_11555 | mul_34_17_n_1077));
 assign mul_34_17_n_4186 = ~((mul_34_17_n_655 & mul_34_17_n_1656) | (mul_34_17_n_2902 & mul_34_17_n_1605));
 assign mul_34_17_n_4185 = ~((mul_34_17_n_667 & mul_34_17_n_644) | (mul_34_17_n_2914 & mul_34_17_n_1248));
 assign mul_34_17_n_4184 = ((mul_34_17_n_678 | mul_34_17_n_884) & (mul_34_17_n_11543 | mul_34_17_n_893));
 assign mul_34_17_n_4183 = ~((mul_34_17_n_675 & mul_34_17_n_989) | (mul_34_17_n_2922 & mul_34_17_n_983));
 assign mul_34_17_n_4182 = ~((mul_34_17_n_671 & mul_34_17_n_1082) | (mul_34_17_n_2918 & mul_34_17_n_1091));
 assign mul_34_17_n_4181 = ((mul_34_17_n_657 & mul_34_17_n_1548) | (mul_34_17_n_2904 & mul_34_17_n_1559));
 assign mul_34_17_n_4179 = ~((mul_34_17_n_661 & mul_34_17_n_1380) | (mul_34_17_n_2908 & mul_34_17_n_1429));
 assign mul_34_17_n_4178 = ((mul_34_17_n_1747 & mul_34_17_n_2028) | (mul_34_17_n_11593 & mul_34_17_n_2100));
 assign mul_34_17_n_4176 = ~((mul_34_17_n_671 & mul_34_17_n_1078) | (mul_34_17_n_2918 & mul_34_17_n_1079));
 assign mul_34_17_n_4175 = ~((mul_34_17_n_1735 & mul_34_17_n_2131) | (mul_34_17_n_2896 & mul_34_17_n_2308));
 assign mul_34_17_n_4174 = ((mul_34_17_n_688 | mul_34_17_n_723) & (mul_34_17_n_11528 | mul_34_17_n_725));
 assign mul_34_17_n_4173 = ~((mul_34_17_n_1743 & mul_34_17_n_2449) | (mul_34_17_n_2882 & mul_34_17_n_1876));
 assign mul_34_17_n_4172 = ~((mul_34_17_n_1757 & mul_34_17_n_1679) | (mul_34_17_n_2900 & mul_34_17_n_1632));
 assign mul_34_17_n_4171 = ~((mul_34_17_n_1747 & mul_34_17_n_1690) | (mul_34_17_n_11593 & mul_34_17_n_2453));
 assign mul_34_17_n_4170 = ~((mul_34_17_n_657 & mul_34_17_n_1526) | (mul_34_17_n_2904 & mul_34_17_n_1550));
 assign mul_34_17_n_4168 = ~((mul_34_17_n_1749 & mul_34_17_n_2672) | (mul_34_17_n_2890 & mul_34_17_n_2101));
 assign mul_34_17_n_4167 = ~((mul_34_17_n_667 & mul_34_17_n_1216) | (mul_34_17_n_2914 & mul_34_17_n_1190));
 assign mul_34_17_n_4166 = ~((mul_34_17_n_687 & mul_34_17_n_650) | (mul_34_17_n_2933 & mul_34_17_n_1337));
 assign mul_34_17_n_4164 = ~((mul_34_17_n_1751 & mul_34_17_n_2654) | (mul_34_17_n_2880 & mul_34_17_n_2669));
 assign mul_34_17_n_4163 = ((mul_34_17_n_1734 | mul_34_17_n_2194) & (mul_34_17_n_11588 | mul_34_17_n_2197));
 assign mul_34_17_n_4162 = ~((mul_34_17_n_677 & mul_34_17_n_928) | (mul_34_17_n_2924 & mul_34_17_n_944));
 assign mul_34_17_n_4161 = ~((mul_34_17_n_1757 & mul_34_17_n_1280) | (mul_34_17_n_2900 & mul_34_17_n_1774));
 assign mul_34_17_n_4160 = ~((mul_34_17_n_687 & mul_34_17_n_712) | (mul_34_17_n_2933 & mul_34_17_n_740));
 assign mul_34_17_n_4159 = ~((mul_34_17_n_665 & mul_34_17_n_1299) | (mul_34_17_n_2912 & mul_34_17_n_1283));
 assign mul_34_17_n_4158 = ~((mul_34_17_n_669 & mul_34_17_n_643) | (mul_34_17_n_2916 & mul_34_17_n_1180));
 assign mul_34_17_n_4157 = ~((mul_34_17_n_677 & mul_34_17_n_943) | (mul_34_17_n_2924 & mul_34_17_n_963));
 assign mul_34_17_n_4156 = ~((mul_34_17_n_1739 & mul_34_17_n_2543) | (mul_34_17_n_2884 & mul_34_17_n_2311));
 assign mul_34_17_n_4155 = ~((mul_34_17_n_677 & mul_34_17_n_639) | (mul_34_17_n_2924 & mul_34_17_n_938));
 assign mul_34_17_n_4154 = ~((mul_34_17_n_1755 & mul_34_17_n_2170) | (mul_34_17_n_2898 & mul_34_17_n_1889));
 assign mul_34_17_n_4152 = ~((mul_34_17_n_525 | mul_34_17_n_529) & (mul_34_17_n_2880 | mul_34_17_n_1751));
 assign mul_34_17_n_4151 = ~((mul_34_17_n_687 & mul_34_17_n_1337) | (mul_34_17_n_2933 & mul_34_17_n_1385));
 assign mul_34_17_n_4150 = ~((mul_34_17_n_665 & mul_34_17_n_1301) | (mul_34_17_n_2912 & mul_34_17_n_1269));
 assign mul_34_17_n_4149 = ((mul_34_17_n_654 | mul_34_17_n_1591) & (mul_34_17_n_11579 | mul_34_17_n_1615));
 assign mul_34_17_n_4148 = ~((mul_34_17_n_669 & mul_34_17_n_1163) | (mul_34_17_n_2916 & mul_34_17_n_1177));
 assign mul_34_17_n_4147 = ((mul_34_17_n_658 | mul_34_17_n_1466) & (mul_34_17_n_11573 | mul_34_17_n_1510));
 assign mul_34_17_n_4146 = ((mul_34_17_n_1744 | mul_34_17_n_1919) & (mul_34_17_n_11600 | mul_34_17_n_2317));
 assign mul_34_17_n_4145 = ~((mul_34_17_n_1751 & mul_34_17_n_2343) | (mul_34_17_n_2880 & mul_34_17_n_2054));
 assign mul_34_17_n_4144 = ~((mul_34_17_n_657 & mul_34_17_n_1561) | (mul_34_17_n_2904 & mul_34_17_n_1558));
 assign mul_34_17_n_4143 = ~((mul_34_17_n_659 & mul_34_17_n_1511) | (mul_34_17_n_2906 & mul_34_17_n_1458));
 assign mul_34_17_n_4142 = ~((mul_34_17_n_659 & mul_34_17_n_1462) | (mul_34_17_n_2906 & mul_34_17_n_1447));
 assign mul_34_17_n_4141 = ((mul_34_17_n_1754 | mul_34_17_n_1884) & (mul_34_17_n_11585 | mul_34_17_n_2420));
 assign mul_34_17_n_4140 = ~((mul_34_17_n_679 & mul_34_17_n_915) | (mul_34_17_n_2926 & mul_34_17_n_916));
 assign mul_34_17_n_4139 = ((mul_34_17_n_682 | mul_34_17_n_818) & (mul_34_17_n_11537 | mul_34_17_n_819));
 assign mul_34_17_n_4138 = ~((mul_34_17_n_523 | mul_34_17_n_526) & (mul_34_17_n_2894 | mul_34_17_n_1737));
 assign mul_34_17_n_4137 = ((mul_34_17_n_1734 | mul_34_17_n_2512) & (mul_34_17_n_11588 | mul_34_17_n_2009));
 assign mul_34_17_n_4136 = ~((mul_34_17_n_527 | mul_34_17_n_528) & (mul_34_17_n_2884 | mul_34_17_n_1739));
 assign mul_34_17_n_4135 = ((mul_34_17_n_1753 & mul_34_17_n_2243) | (mul_34_17_n_2878 & mul_34_17_n_2092));
 assign mul_34_17_n_4134 = ((mul_34_17_n_655 & mul_34_17_n_1633) | (mul_34_17_n_2902 & mul_34_17_n_1610));
 assign mul_34_17_n_4132 = ~((mul_34_17_n_667 & mul_34_17_n_1240) | (mul_34_17_n_2914 & mul_34_17_n_1245));
 assign mul_34_17_n_4131 = ~((mul_34_17_n_1751 & mul_34_17_n_2180) | (mul_34_17_n_2880 & mul_34_17_n_2036));
 assign mul_34_17_n_4130 = ~((mul_34_17_n_659 & mul_34_17_n_1494) | (mul_34_17_n_2906 & mul_34_17_n_1513));
 assign mul_34_17_n_4129 = ~((mul_34_17_n_673 & mul_34_17_n_1025) | (mul_34_17_n_2920 & mul_34_17_n_1036));
 assign mul_34_17_n_4128 = ~((mul_34_17_n_1739 & mul_34_17_n_2579) | (mul_34_17_n_2884 & mul_34_17_n_1847));
 assign mul_34_17_n_4127 = ~((mul_34_17_n_663 & mul_34_17_n_1310) | (mul_34_17_n_2910 & mul_34_17_n_1311));
 assign mul_34_17_n_4126 = ((mul_34_17_n_1736 | mul_34_17_n_1940) & (mul_34_17_n_11591 | mul_34_17_n_1976));
 assign mul_34_17_n_4125 = ~((mul_34_17_n_661 & mul_34_17_n_1383) | (mul_34_17_n_2908 & mul_34_17_n_1427));
 assign mul_34_17_n_4124 = ((mul_34_17_n_662 | mul_34_17_n_1341) & (mul_34_17_n_11567 | mul_34_17_n_1314));
 assign mul_34_17_n_4123 = ~((mul_34_17_n_671 & mul_34_17_n_1107) | (mul_34_17_n_2918 & mul_34_17_n_1080));
 assign mul_34_17_n_4122 = ~((mul_34_17_n_659 & mul_34_17_n_1458) | (mul_34_17_n_2906 & mul_34_17_n_1452));
 assign mul_34_17_n_4121 = ~((mul_34_17_n_1757 & mul_34_17_n_2257) | (mul_34_17_n_2900 & mul_34_17_n_1764));
 assign mul_34_17_n_4120 = ((mul_34_17_n_686 | mul_34_17_n_733) & (mul_34_17_n_11531 | mul_34_17_n_716));
 assign mul_34_17_n_4119 = ((mul_34_17_n_1753 & mul_34_17_n_2008) | (mul_34_17_n_2878 & mul_34_17_n_2260));
 assign mul_34_17_n_4118 = ~((mul_34_17_n_677 & mul_34_17_n_930) | (mul_34_17_n_2924 & mul_34_17_n_937));
 assign mul_34_17_n_4117 = ((mul_34_17_n_660 | mul_34_17_n_1444) & (mul_34_17_n_11570 | mul_34_17_n_1432));
 assign mul_34_17_n_4116 = ((mul_34_17_n_661 & mul_34_17_n_1441) | (mul_34_17_n_2908 & mul_34_17_n_1404));
 assign mul_34_17_n_4115 = ~((mul_34_17_n_1753 & mul_34_17_n_2319) | (mul_34_17_n_2878 & mul_34_17_n_2008));
 assign mul_34_17_n_4114 = ((mul_34_17_n_1750 | mul_34_17_n_2413) & (mul_34_17_n_11612 | mul_34_17_n_1907));
 assign mul_34_17_n_4113 = ((mul_34_17_n_1754 | mul_34_17_n_2090) & (mul_34_17_n_11585 | mul_34_17_n_2495));
 assign mul_34_17_n_4112 = ((mul_34_17_n_491 & mul_34_17_n_490) | (mul_34_17_n_11597 & mul_34_17_n_1748));
 assign mul_34_17_n_4111 = ~((mul_34_17_n_1741 & mul_34_17_n_2476) | (mul_34_17_n_2886 & mul_34_17_n_2363));
 assign mul_34_17_n_4109 = ((mul_34_17_n_682 | mul_34_17_n_805) & (mul_34_17_n_11537 | mul_34_17_n_825));
 assign mul_34_17_n_4108 = ((mul_34_17_n_654 | mul_34_17_n_1609) & (mul_34_17_n_11579 | mul_34_17_n_1607));
 assign mul_34_17_n_4107 = ((mul_34_17_n_1735 & mul_34_17_n_1693) | (mul_34_17_n_2896 & mul_34_17_n_2694));
 assign mul_34_17_n_4106 = ~((mul_34_17_n_667 & mul_34_17_n_1247) | (mul_34_17_n_2914 & mul_34_17_n_1189));
 assign mul_34_17_n_4105 = ((mul_34_17_n_1743 & mul_34_17_n_2118) | (mul_34_17_n_2882 & mul_34_17_n_2282));
 assign mul_34_17_n_4104 = ~((mul_34_17_n_655 & mul_34_17_n_1637) | (mul_34_17_n_2902 & mul_34_17_n_1654));
 assign mul_34_17_n_4103 = ((mul_34_17_n_1753 & mul_34_17_n_1877) | (mul_34_17_n_2878 & mul_34_17_n_2428));
 assign mul_34_17_n_4102 = ((mul_34_17_n_667 & mul_34_17_n_1248) | (mul_34_17_n_2914 & mul_34_17_n_1204));
 assign mul_34_17_n_4100 = ((mul_34_17_n_519 & mul_34_17_n_521) | (mul_34_17_n_11653 & mul_34_17_n_1746));
 assign mul_34_17_n_4099 = ~((mul_34_17_n_679 & mul_34_17_n_901) | (mul_34_17_n_2926 & mul_34_17_n_907));
 assign mul_34_17_n_4098 = ~((mul_34_17_n_665 & mul_34_17_n_1289) | (mul_34_17_n_2912 & mul_34_17_n_1253));
 assign mul_34_17_n_4096 = ~((mul_34_17_n_1741 & mul_34_17_n_1947) | (mul_34_17_n_2886 & mul_34_17_n_2418));
 assign mul_34_17_n_4095 = ~((mul_34_17_n_671 & mul_34_17_n_1093) | (mul_34_17_n_2918 & mul_34_17_n_1082));
 assign mul_34_17_n_4094 = ~((mul_34_17_n_663 & mul_34_17_n_646) | (mul_34_17_n_2910 & mul_34_17_n_1328));
 assign mul_34_17_n_4093 = ((mul_34_17_n_656 | mul_34_17_n_1545) & (mul_34_17_n_11576 | mul_34_17_n_1530));
 assign mul_34_17_n_4092 = ((mul_34_17_n_680 | mul_34_17_n_836) & (mul_34_17_n_11540 | mul_34_17_n_851));
 assign mul_34_17_n_4091 = ((mul_34_17_n_676 | mul_34_17_n_964) & (mul_34_17_n_11546 | mul_34_17_n_949));
 assign mul_34_17_n_4090 = ~((mul_34_17_n_669 & mul_34_17_n_1166) | (mul_34_17_n_2916 & mul_34_17_n_1158));
 assign mul_34_17_n_4089 = ((mul_34_17_n_1752 | mul_34_17_n_2402) & (mul_34_17_n_11615 | mul_34_17_n_2401));
 assign mul_34_17_n_4088 = ((mul_34_17_n_1737 & mul_34_17_n_2056) | (mul_34_17_n_2894 & mul_34_17_n_2653));
 assign mul_34_17_n_4087 = ~((mul_34_17_n_657 & mul_34_17_n_649) | (mul_34_17_n_2904 & mul_34_17_n_1583));
 assign mul_34_17_n_4086 = ~((mul_34_17_n_1757 & mul_34_17_n_1776) | (mul_34_17_n_2900 & mul_34_17_n_1763));
 assign mul_34_17_n_4085 = ((mul_34_17_n_663 & mul_34_17_n_1352) | (mul_34_17_n_2910 & mul_34_17_n_1340));
 assign mul_34_17_n_4084 = ((mul_34_17_n_1747 & mul_34_17_n_1931) | (mul_34_17_n_11593 & mul_34_17_n_2276));
 assign mul_34_17_n_4083 = ((mul_34_17_n_682 | mul_34_17_n_833) & (mul_34_17_n_11537 | mul_34_17_n_821));
 assign mul_34_17_n_4082 = ((mul_34_17_n_658 | mul_34_17_n_1451) & (mul_34_17_n_11573 | mul_34_17_n_1493));
 assign mul_34_17_n_4081 = ((mul_34_17_n_489 | mul_34_17_n_488) & (mul_34_17_n_2888 | mul_34_17_n_1745));
 assign mul_34_17_n_4080 = ~((mul_34_17_n_691 & mul_34_17_n_634) | (mul_34_17_n_2936 & mul_34_17_n_693));
 assign mul_34_17_n_4079 = ((mul_34_17_n_662 | mul_34_17_n_1347) & (mul_34_17_n_11567 | mul_34_17_n_1341));
 assign mul_34_17_n_4078 = ~((mul_34_17_n_677 & mul_34_17_n_952) | (mul_34_17_n_2924 & mul_34_17_n_939));
 assign mul_34_17_n_4077 = ((mul_34_17_n_664 | mul_34_17_n_1281) & (mul_34_17_n_11564 | mul_34_17_n_1250));
 assign mul_34_17_n_4076 = ((mul_34_17_n_520 & mul_34_17_n_530) | (mul_34_17_n_11588 & mul_34_17_n_1734));
 assign mul_34_17_n_4075 = ~((mul_34_17_n_1749 & mul_34_17_n_2576) | (mul_34_17_n_2890 & mul_34_17_n_2143));
 assign mul_34_17_n_4074 = ((mul_34_17_n_1752 | mul_34_17_n_2401) & (mul_34_17_n_11615 | mul_34_17_n_2619));
 assign mul_34_17_n_4073 = ~((mul_34_17_n_691 & mul_34_17_n_1058) | (mul_34_17_n_2936 & mul_34_17_n_751));
 assign mul_34_17_n_4071 = ~((mul_34_17_n_1737 & mul_34_17_n_1962) | (mul_34_17_n_2894 & mul_34_17_n_1866));
 assign mul_34_17_n_4070 = ~((mul_34_17_n_1755 & mul_34_17_n_2676) | (mul_34_17_n_2898 & mul_34_17_n_2547));
 assign mul_34_17_n_4069 = ((mul_34_17_n_1740 | mul_34_17_n_2386) & (mul_34_17_n_11603 | mul_34_17_n_1923));
 assign mul_34_17_n_4067 = ~((mul_34_17_n_1749 & mul_34_17_n_2415) | (mul_34_17_n_2890 & mul_34_17_n_2235));
 assign mul_34_17_n_4066 = ~((mul_34_17_n_1741 & mul_34_17_n_2120) | (mul_34_17_n_2886 & mul_34_17_n_2279));
 assign mul_34_17_n_4065 = ((mul_34_17_n_655 & mul_34_17_n_1664) | (mul_34_17_n_2902 & mul_34_17_n_1663));
 assign mul_34_17_n_4064 = ~((mul_34_17_n_671 & mul_34_17_n_1086) | (mul_34_17_n_2918 & mul_34_17_n_1116));
 assign mul_34_17_n_4063 = ((mul_34_17_n_675 & mul_34_17_n_1010) | (mul_34_17_n_2922 & mul_34_17_n_994));
 assign mul_34_17_n_4062 = ((mul_34_17_n_657 & mul_34_17_n_1567) | (mul_34_17_n_2904 & mul_34_17_n_1526));
 assign mul_34_17_n_4061 = ~((mul_34_17_n_657 & mul_34_17_n_1569) | (mul_34_17_n_2904 & mul_34_17_n_1571));
 assign mul_34_17_n_4060 = ~((mul_34_17_n_659 & mul_34_17_n_1514) | (mul_34_17_n_2906 & mul_34_17_n_1459));
 assign mul_34_17_n_4059 = ~((mul_34_17_n_677 & mul_34_17_n_923) | (mul_34_17_n_2924 & mul_34_17_n_925));
 assign mul_34_17_n_4058 = ~((mul_34_17_n_681 & mul_34_17_n_855) | (mul_34_17_n_2928 & mul_34_17_n_839));
 assign mul_34_17_n_4057 = ((mul_34_17_n_1757 & mul_34_17_n_1683) | (mul_34_17_n_2900 & mul_34_17_n_1959));
 assign mul_34_17_n_4056 = ~((mul_34_17_n_665 & mul_34_17_n_1292) | (mul_34_17_n_2912 & mul_34_17_n_1290));
 assign mul_34_17_n_4055 = ~((mul_34_17_n_657 & mul_34_17_n_1574) | (mul_34_17_n_2904 & mul_34_17_n_1541));
 assign mul_34_17_n_4054 = ~((mul_34_17_n_1749 & mul_34_17_n_2665) | (mul_34_17_n_2890 & mul_34_17_n_1930));
 assign mul_34_17_n_4053 = ~((mul_34_17_n_1743 & mul_34_17_n_2301) | (mul_34_17_n_2882 & mul_34_17_n_2240));
 assign mul_34_17_n_4052 = ~((mul_34_17_n_1757 & mul_34_17_n_1680) | (mul_34_17_n_2900 & mul_34_17_n_1776));
 assign mul_34_17_n_4051 = ((mul_34_17_n_691 & mul_34_17_n_732) | (mul_34_17_n_2936 & mul_34_17_n_720));
 assign mul_34_17_n_4050 = ~((mul_34_17_n_691 & mul_34_17_n_710) | (mul_34_17_n_2936 & mul_34_17_n_721));
 assign mul_34_17_n_4049 = ~(mul_34_17_n_2740 ^ mul_34_17_n_2855);
 assign mul_34_17_n_4048 = ~((mul_34_17_n_492 | mul_34_17_n_487) & (mul_34_17_n_2882 | mul_34_17_n_1743));
 assign mul_34_17_n_4047 = ~((mul_34_17_n_1749 & mul_34_17_n_2534) | (mul_34_17_n_2890 & mul_34_17_n_2369));
 assign mul_34_17_n_4046 = ~((mul_34_17_n_685 & mul_34_17_n_796) | (mul_34_17_n_2931 & mul_34_17_n_792));
 assign mul_34_17_n_4044 = ((mul_34_17_n_1736 | mul_34_17_n_2332) & (mul_34_17_n_11591 | mul_34_17_n_2269));
 assign mul_34_17_n_4043 = ~((mul_34_17_n_1755 & mul_34_17_n_2667) | (mul_34_17_n_2898 & mul_34_17_n_2255));
 assign mul_34_17_n_4042 = ~((mul_34_17_n_522 | mul_34_17_n_524) & (mul_34_17_n_2886 | mul_34_17_n_1741));
 assign mul_34_17_n_4041 = ~((mul_34_17_n_659 & mul_34_17_n_1452) | (mul_34_17_n_2906 & mul_34_17_n_1506));
 assign mul_34_17_n_4040 = ~((mul_34_17_n_671 & mul_34_17_n_1104) | (mul_34_17_n_2918 & mul_34_17_n_1067));
 assign mul_34_17_n_4039 = ~((mul_34_17_n_667 & mul_34_17_n_1214) | (mul_34_17_n_2914 & mul_34_17_n_1187));
 assign mul_34_17_n_4038 = ((mul_34_17_n_1736 | mul_34_17_n_2347) & (mul_34_17_n_11591 | mul_34_17_n_2380));
 assign mul_34_17_n_4037 = ((mul_34_17_n_658 | mul_34_17_n_1501) & (mul_34_17_n_11573 | mul_34_17_n_1478));
 assign mul_34_17_n_4036 = ~((mul_34_17_n_669 & mul_34_17_n_1138) | (mul_34_17_n_2916 & mul_34_17_n_1155));
 assign mul_34_17_n_4034 = ((mul_34_17_n_662 | mul_34_17_n_1333) & (mul_34_17_n_11567 | mul_34_17_n_1347));
 assign mul_34_17_n_4033 = ~((mul_34_17_n_675 & mul_34_17_n_996) | (mul_34_17_n_2922 & mul_34_17_n_1000));
 assign mul_34_17_n_4032 = ~((mul_34_17_n_1741 & mul_34_17_n_2541) | (mul_34_17_n_2886 & mul_34_17_n_2589));
 assign mul_34_17_n_4031 = ~((mul_34_17_n_1749 & mul_34_17_n_2604) | (mul_34_17_n_2890 & mul_34_17_n_2432));
 assign mul_34_17_n_4030 = ((mul_34_17_n_1756 | mul_34_17_n_1686) & (mul_34_17_n_11582 | mul_34_17_n_2377));
 assign mul_34_17_n_4029 = ((mul_34_17_n_682 | mul_34_17_n_823) & (mul_34_17_n_11537 | mul_34_17_n_818));
 assign mul_34_17_n_4028 = ~((mul_34_17_n_1755 & mul_34_17_n_2059) | (mul_34_17_n_2898 & mul_34_17_n_2148));
 assign mul_34_17_n_4027 = ~((mul_34_17_n_679 & mul_34_17_n_889) | (mul_34_17_n_2926 & mul_34_17_n_898));
 assign mul_34_17_n_4026 = ((mul_34_17_n_1736 | mul_34_17_n_2178) & (mul_34_17_n_11591 | mul_34_17_n_2376));
 assign mul_34_17_n_4025 = ((mul_34_17_n_684 | mul_34_17_n_766) & (mul_34_17_n_11534 | mul_34_17_n_791));
 assign mul_34_17_n_4023 = ((mul_34_17_n_664 | mul_34_17_n_1307) & (mul_34_17_n_11564 | mul_34_17_n_1285));
 assign mul_34_17_n_4022 = ((mul_34_17_n_686 | mul_34_17_n_713) & (mul_34_17_n_11531 | mul_34_17_n_733));
 assign mul_34_17_n_4021 = ~(mul_34_17_n_2999 | mul_34_17_n_2749);
 assign mul_34_17_n_4020 = ~((mul_34_17_n_1747 & mul_34_17_n_2108) | (mul_34_17_n_11593 & mul_34_17_n_2617));
 assign mul_34_17_n_4019 = ~((mul_34_17_n_1757 & mul_34_17_n_1764) | (mul_34_17_n_2900 & mul_34_17_n_1771));
 assign mul_34_17_n_4017 = ~((mul_34_17_n_1755 & mul_34_17_n_2027) | (mul_34_17_n_2898 & mul_34_17_n_2667));
 assign mul_34_17_n_4015 = ((mul_34_17_n_1738 | mul_34_17_n_1996) & (mul_34_17_n_11606 | mul_34_17_n_2327));
 assign mul_34_17_n_4013 = ~((mul_34_17_n_1747 & mul_34_17_n_2174) | (mul_34_17_n_11593 & mul_34_17_n_2562));
 assign mul_34_17_n_4011 = ((mul_34_17_n_1738 | mul_34_17_n_2487) & (mul_34_17_n_11606 | mul_34_17_n_2105));
 assign mul_34_17_n_4010 = ~((mul_34_17_n_657 & mul_34_17_n_1543) | (mul_34_17_n_2904 & mul_34_17_n_1552));
 assign mul_34_17_n_4009 = ((mul_34_17_n_1742 | mul_34_17_n_2058) & (mul_34_17_n_11609 | mul_34_17_n_2408));
 assign mul_34_17_n_4008 = ~((mul_34_17_n_1739 & mul_34_17_n_2389) | (mul_34_17_n_2884 & mul_34_17_n_2390));
 assign mul_34_17_n_4006 = ((mul_34_17_n_1740 | mul_34_17_n_2057) & (mul_34_17_n_11603 | mul_34_17_n_2386));
 assign mul_34_17_n_4004 = ((mul_34_17_n_670 | mul_34_17_n_1115) & (mul_34_17_n_11555 | mul_34_17_n_1069));
 assign mul_34_17_n_4003 = ~((mul_34_17_n_1752 | mul_34_17_n_2107) & (mul_34_17_n_11615 | mul_34_17_n_2402));
 assign mul_34_17_n_4002 = ~((mul_34_17_n_669 & mul_34_17_n_1180) | (mul_34_17_n_2916 & mul_34_17_n_1144));
 assign mul_34_17_n_4001 = ~((mul_34_17_n_1739 & mul_34_17_n_1841) | (mul_34_17_n_2884 & mul_34_17_n_2344));
 assign mul_34_17_n_3999 = ~((mul_34_17_n_677 & mul_34_17_n_966) | (mul_34_17_n_2924 & mul_34_17_n_948));
 assign mul_34_17_n_3998 = ~((mul_34_17_n_1745 & mul_34_17_n_2530) | (mul_34_17_n_2888 & mul_34_17_n_1875));
 assign mul_34_17_n_3996 = ((mul_34_17_n_668 | mul_34_17_n_1171) & (mul_34_17_n_11558 | mul_34_17_n_1174));
 assign mul_34_17_n_3994 = ((mul_34_17_n_678 | mul_34_17_n_917) & (mul_34_17_n_11543 | mul_34_17_n_900));
 assign mul_34_17_n_3993 = ~((mul_34_17_n_1737 & mul_34_17_n_2270) | (mul_34_17_n_2894 & mul_34_17_n_2618));
 assign mul_34_17_n_3992 = ~((mul_34_17_n_1745 & mul_34_17_n_2518) | (mul_34_17_n_2888 & mul_34_17_n_2303));
 assign mul_34_17_n_3991 = ~((mul_34_17_n_1757 & mul_34_17_n_1763) | (mul_34_17_n_2900 & mul_34_17_n_1666));
 assign mul_34_17_n_3990 = ~((mul_34_17_n_1747 & mul_34_17_n_1945) | (mul_34_17_n_11593 & mul_34_17_n_2647));
 assign mul_34_17_n_3988 = ((mul_34_17_n_674 | mul_34_17_n_1013) & (mul_34_17_n_11549 | mul_34_17_n_984));
 assign mul_34_17_n_3987 = ~((mul_34_17_n_1737 & mul_34_17_n_2251) | (mul_34_17_n_2894 & mul_34_17_n_2411));
 assign mul_34_17_n_3986 = ~((mul_34_17_n_1751 & mul_34_17_n_2054) | (mul_34_17_n_2880 & mul_34_17_n_2644));
 assign mul_34_17_n_3983 = ~((mul_34_17_n_1749 & mul_34_17_n_1930) | (mul_34_17_n_2890 & mul_34_17_n_2507));
 assign mul_34_17_n_3981 = ((mul_34_17_n_1742 | mul_34_17_n_2371) & (mul_34_17_n_11609 | mul_34_17_n_1943));
 assign mul_34_17_n_3980 = ((mul_34_17_n_666 | mul_34_17_n_1239) & (mul_34_17_n_11561 | mul_34_17_n_1230));
 assign mul_34_17_n_3979 = ~(mul_34_17_n_2869 ^ mul_34_17_n_2955);
 assign mul_34_17_n_3978 = ~((mul_34_17_n_675 & mul_34_17_n_994) | (mul_34_17_n_2922 & mul_34_17_n_1002));
 assign mul_34_17_n_3977 = ~((mul_34_17_n_1755 & mul_34_17_n_2255) | (mul_34_17_n_2898 & mul_34_17_n_1849));
 assign mul_34_17_n_3976 = ~((mul_34_17_n_1749 & mul_34_17_n_2196) | (mul_34_17_n_2890 & mul_34_17_n_1994));
 assign mul_34_17_n_3975 = ~((mul_34_17_n_677 & mul_34_17_n_961) | (mul_34_17_n_2924 & mul_34_17_n_951));
 assign mul_34_17_n_3974 = ((mul_34_17_n_1757 & mul_34_17_n_1674) | (mul_34_17_n_2900 & mul_34_17_n_799));
 assign mul_34_17_n_3973 = ~(mul_34_17_n_2947 ^ mul_34_17_n_2859);
 assign mul_34_17_n_3972 = ~((mul_34_17_n_679 & mul_34_17_n_880) | (mul_34_17_n_2926 & mul_34_17_n_905));
 assign mul_34_17_n_3971 = ((mul_34_17_n_1753 & mul_34_17_n_2137) | (mul_34_17_n_2878 & mul_34_17_n_1995));
 assign mul_34_17_n_3970 = ((mul_34_17_n_671 & mul_34_17_n_1080) | (mul_34_17_n_2918 & mul_34_17_n_1089));
 assign mul_34_17_n_3969 = ~((mul_34_17_n_1747 & mul_34_17_n_2226) | (mul_34_17_n_11593 & mul_34_17_n_1990));
 assign mul_34_17_n_3967 = ~((mul_34_17_n_1747 & mul_34_17_n_2404) | (mul_34_17_n_11593 & mul_34_17_n_2288));
 assign mul_34_17_n_3966 = ~((mul_34_17_n_1743 & mul_34_17_n_1871) | (mul_34_17_n_2882 & mul_34_17_n_2664));
 assign mul_34_17_n_3964 = ~((mul_34_17_n_691 & mul_34_17_n_699) | (mul_34_17_n_2936 & mul_34_17_n_734));
 assign mul_34_17_n_3962 = ~((mul_34_17_n_1741 & mul_34_17_n_1989) | (mul_34_17_n_2886 & mul_34_17_n_2473));
 assign mul_34_17_n_3961 = ~((mul_34_17_n_673 & mul_34_17_n_1061) | (mul_34_17_n_2920 & mul_34_17_n_1055));
 assign mul_34_17_n_3942 = ~mul_34_17_n_3941;
 assign mul_34_17_n_3940 = ~mul_34_17_n_3939;
 assign mul_34_17_n_3921 = ~mul_34_17_n_3920;
 assign mul_34_17_n_3918 = ~mul_34_17_n_3917;
 assign mul_34_17_n_3905 = ~mul_34_17_n_3904;
 assign mul_34_17_n_3901 = ~mul_34_17_n_3900;
 assign mul_34_17_n_3897 = ~mul_34_17_n_3896;
 assign mul_34_17_n_3890 = ~mul_34_17_n_3889;
 assign mul_34_17_n_3863 = ~mul_34_17_n_3862;
 assign mul_34_17_n_3860 = ~mul_34_17_n_3859;
 assign mul_34_17_n_3857 = ~mul_34_17_n_3856;
 assign mul_34_17_n_3851 = ~mul_34_17_n_3850;
 assign mul_34_17_n_3849 = ~mul_34_17_n_3848;
 assign mul_34_17_n_3846 = ~mul_34_17_n_3845;
 assign mul_34_17_n_3838 = ~mul_34_17_n_3837;
 assign mul_34_17_n_3823 = ~mul_34_17_n_3822;
 assign mul_34_17_n_3820 = ~mul_34_17_n_3819;
 assign mul_34_17_n_3805 = ~mul_34_17_n_3804;
 assign mul_34_17_n_3803 = ~mul_34_17_n_3802;
 assign mul_34_17_n_3780 = ~mul_34_17_n_3779;
 assign mul_34_17_n_3777 = ~mul_34_17_n_3776;
 assign mul_34_17_n_3773 = ~mul_34_17_n_3772;
 assign mul_34_17_n_3767 = ~mul_34_17_n_3766;
 assign mul_34_17_n_3763 = ~mul_34_17_n_3762;
 assign mul_34_17_n_3745 = ~mul_34_17_n_3744;
 assign mul_34_17_n_3722 = ~mul_34_17_n_3721;
 assign mul_34_17_n_3702 = ~mul_34_17_n_3701;
 assign mul_34_17_n_3697 = ~mul_34_17_n_3696;
 assign mul_34_17_n_3695 = ~mul_34_17_n_3694;
 assign mul_34_17_n_3688 = ~mul_34_17_n_3687;
 assign mul_34_17_n_3686 = ~mul_34_17_n_3685;
 assign mul_34_17_n_3683 = ~mul_34_17_n_3682;
 assign mul_34_17_n_3680 = ~mul_34_17_n_3679;
 assign mul_34_17_n_3670 = ~mul_34_17_n_3669;
 assign mul_34_17_n_3663 = ~mul_34_17_n_3662;
 assign mul_34_17_n_3644 = ~mul_34_17_n_3643;
 assign mul_34_17_n_3636 = ~mul_34_17_n_3635;
 assign mul_34_17_n_3631 = ~mul_34_17_n_3630;
 assign mul_34_17_n_3627 = ~mul_34_17_n_3626;
 assign mul_34_17_n_3615 = ~mul_34_17_n_3614;
 assign mul_34_17_n_3613 = ~mul_34_17_n_3612;
 assign mul_34_17_n_3604 = ~mul_34_17_n_3603;
 assign mul_34_17_n_3596 = ~mul_34_17_n_3595;
 assign mul_34_17_n_3593 = ~mul_34_17_n_3592;
 assign mul_34_17_n_3591 = ~mul_34_17_n_3590;
 assign mul_34_17_n_3589 = ~mul_34_17_n_3588;
 assign mul_34_17_n_3577 = ~mul_34_17_n_3576;
 assign mul_34_17_n_3569 = ~mul_34_17_n_3568;
 assign mul_34_17_n_3557 = ~mul_34_17_n_3556;
 assign mul_34_17_n_3555 = ~mul_34_17_n_3554;
 assign mul_34_17_n_3552 = ~mul_34_17_n_3551;
 assign mul_34_17_n_3545 = ~mul_34_17_n_3544;
 assign mul_34_17_n_3543 = ~mul_34_17_n_3542;
 assign mul_34_17_n_3540 = ~mul_34_17_n_3539;
 assign mul_34_17_n_3535 = ~mul_34_17_n_3534;
 assign mul_34_17_n_3532 = ~mul_34_17_n_3531;
 assign mul_34_17_n_3528 = ~mul_34_17_n_3527;
 assign mul_34_17_n_3524 = ~mul_34_17_n_3523;
 assign mul_34_17_n_3514 = ~mul_34_17_n_3513;
 assign mul_34_17_n_3504 = ~mul_34_17_n_3503;
 assign mul_34_17_n_3502 = ~mul_34_17_n_3501;
 assign mul_34_17_n_3498 = ~mul_34_17_n_3497;
 assign mul_34_17_n_3495 = ~mul_34_17_n_3494;
 assign mul_34_17_n_3443 = ~mul_34_17_n_3442;
 assign mul_34_17_n_3416 = ~mul_34_17_n_3415;
 assign mul_34_17_n_3404 = ~mul_34_17_n_3403;
 assign mul_34_17_n_3400 = ~mul_34_17_n_3399;
 assign mul_34_17_n_3398 = ~mul_34_17_n_3397;
 assign mul_34_17_n_3396 = ~mul_34_17_n_3395;
 assign mul_34_17_n_3394 = ~mul_34_17_n_3393;
 assign mul_34_17_n_3392 = ~mul_34_17_n_3391;
 assign mul_34_17_n_3390 = ~mul_34_17_n_3389;
 assign mul_34_17_n_3388 = ~mul_34_17_n_3387;
 assign mul_34_17_n_3369 = ~mul_34_17_n_3368;
 assign mul_34_17_n_3352 = ~mul_34_17_n_3351;
 assign mul_34_17_n_3350 = ~mul_34_17_n_3349;
 assign mul_34_17_n_3342 = ~mul_34_17_n_3341;
 assign mul_34_17_n_3337 = ~mul_34_17_n_3336;
 assign mul_34_17_n_3331 = ~mul_34_17_n_3330;
 assign mul_34_17_n_3325 = ~mul_34_17_n_3324;
 assign mul_34_17_n_3318 = ~mul_34_17_n_3317;
 assign mul_34_17_n_3312 = ~mul_34_17_n_3311;
 assign mul_34_17_n_3292 = ~mul_34_17_n_3291;
 assign mul_34_17_n_3290 = ~mul_34_17_n_3289;
 assign mul_34_17_n_3272 = ~mul_34_17_n_3271;
 assign mul_34_17_n_3270 = ~mul_34_17_n_3269;
 assign mul_34_17_n_3268 = ~mul_34_17_n_3267;
 assign mul_34_17_n_3260 = ~mul_34_17_n_3259;
 assign mul_34_17_n_3247 = ~mul_34_17_n_3246;
 assign mul_34_17_n_3245 = ~mul_34_17_n_3244;
 assign mul_34_17_n_3242 = ~mul_34_17_n_3241;
 assign mul_34_17_n_3240 = ~mul_34_17_n_3239;
 assign mul_34_17_n_3237 = ~mul_34_17_n_3236;
 assign mul_34_17_n_3229 = ~mul_34_17_n_3228;
 assign mul_34_17_n_3208 = ~mul_34_17_n_3207;
 assign mul_34_17_n_3203 = ~mul_34_17_n_3202;
 assign mul_34_17_n_3201 = ~mul_34_17_n_3200;
 assign mul_34_17_n_3199 = ~mul_34_17_n_3198;
 assign mul_34_17_n_3196 = ~mul_34_17_n_3195;
 assign mul_34_17_n_3181 = ~mul_34_17_n_3180;
 assign mul_34_17_n_3167 = ~mul_34_17_n_3166;
 assign mul_34_17_n_3165 = ~mul_34_17_n_3164;
 assign mul_34_17_n_3163 = ~mul_34_17_n_3162;
 assign mul_34_17_n_3161 = ~mul_34_17_n_3160;
 assign mul_34_17_n_3153 = ~mul_34_17_n_3152;
 assign mul_34_17_n_3146 = ~mul_34_17_n_3145;
 assign mul_34_17_n_3144 = ~mul_34_17_n_3143;
 assign mul_34_17_n_3142 = ~mul_34_17_n_3141;
 assign mul_34_17_n_3138 = ~mul_34_17_n_3137;
 assign mul_34_17_n_3136 = ~mul_34_17_n_3135;
 assign mul_34_17_n_3133 = ~mul_34_17_n_3132;
 assign mul_34_17_n_3131 = ~mul_34_17_n_3130;
 assign mul_34_17_n_3129 = ~mul_34_17_n_3128;
 assign mul_34_17_n_3116 = ~mul_34_17_n_3115;
 assign mul_34_17_n_3114 = ~mul_34_17_n_3113;
 assign mul_34_17_n_3110 = ~mul_34_17_n_3109;
 assign mul_34_17_n_3100 = ~mul_34_17_n_3099;
 assign mul_34_17_n_3095 = ~mul_34_17_n_3094;
 assign mul_34_17_n_3090 = ~mul_34_17_n_3089;
 assign mul_34_17_n_3081 = ~mul_34_17_n_3080;
 assign mul_34_17_n_3077 = ~mul_34_17_n_3076;
 assign mul_34_17_n_3073 = ~mul_34_17_n_3072;
 assign mul_34_17_n_3071 = ~mul_34_17_n_3070;
 assign mul_34_17_n_3067 = ~mul_34_17_n_3068;
 assign mul_34_17_n_3066 = ~mul_34_17_n_3065;
 assign mul_34_17_n_3064 = ~mul_34_17_n_3063;
 assign mul_34_17_n_3060 = ~mul_34_17_n_3061;
 assign mul_34_17_n_3944 = ~((mul_34_17_n_1749 & mul_34_17_n_2493) | (mul_34_17_n_2890 & mul_34_17_n_1846));
 assign mul_34_17_n_3052 = ~(mul_34_17_n_2714 ^ mul_34_17_n_2841);
 assign mul_34_17_n_3943 = ~((mul_34_17_n_684 | mul_34_17_n_780) & (mul_34_17_n_11534 | mul_34_17_n_778));
 assign mul_34_17_n_3051 = ~((mul_34_17_n_665 & mul_34_17_n_645) | (mul_34_17_n_2912 & mul_34_17_n_1272));
 assign mul_34_17_n_3050 = (mul_34_17_n_2715 ^ mul_34_17_n_2845);
 assign mul_34_17_n_3049 = ((mul_34_17_n_654 | mul_34_17_n_651) & (mul_34_17_n_11579 | mul_34_17_n_1621));
 assign mul_34_17_n_3941 = ((mul_34_17_n_678 | mul_34_17_n_908) & (mul_34_17_n_11543 | mul_34_17_n_876));
 assign mul_34_17_n_3048 = ~(mul_34_17_n_2713 ^ mul_34_17_n_2839);
 assign mul_34_17_n_3939 = ((mul_34_17_n_1750 | mul_34_17_n_2598) & (mul_34_17_n_11612 | mul_34_17_n_2362));
 assign mul_34_17_n_3938 = ((mul_34_17_n_1746 | mul_34_17_n_2560) & (mul_34_17_n_11645 | mul_34_17_n_2081));
 assign mul_34_17_n_3937 = (mul_34_17_n_2741 ^ mul_34_17_n_2821);
 assign mul_34_17_n_3047 = ~(mul_34_17_n_2737 ^ mul_34_17_n_2831);
 assign mul_34_17_n_3936 = ((mul_34_17_n_1744 | mul_34_17_n_2403) & (mul_34_17_n_11600 | mul_34_17_n_2103));
 assign mul_34_17_n_3046 = ~((mul_34_17_n_1757 & mul_34_17_n_653) | (mul_34_17_n_2900 & mul_34_17_n_1680));
 assign mul_34_17_n_3045 = ~(mul_34_17_n_2719 ^ mul_34_17_n_2833);
 assign mul_34_17_n_3935 = ~((mul_34_17_n_1745 & mul_34_17_n_2135) | (mul_34_17_n_2888 & mul_34_17_n_2475));
 assign mul_34_17_n_3044 = (mul_34_17_n_2844 ^ mul_34_17_n_2722);
 assign mul_34_17_n_3934 = (mul_34_17_n_2716 ^ mul_34_17_n_2854);
 assign mul_34_17_n_3933 = ~((mul_34_17_n_1745 & mul_34_17_n_2205) | (mul_34_17_n_2888 & mul_34_17_n_2643));
 assign mul_34_17_n_3932 = ~((mul_34_17_n_691 & mul_34_17_n_693) | (mul_34_17_n_2936 & mul_34_17_n_715));
 assign mul_34_17_n_3931 = ~((mul_34_17_n_690 | mul_34_17_n_702) & (mul_34_17_n_11525 | mul_34_17_n_737));
 assign mul_34_17_n_3043 = (mul_34_17_n_2731 ^ mul_34_17_n_2824);
 assign mul_34_17_n_3930 = ~((mul_34_17_n_1734 | mul_34_17_n_2510) & (mul_34_17_n_11588 | mul_34_17_n_1918));
 assign mul_34_17_n_3929 = ((mul_34_17_n_1744 | mul_34_17_n_2015) & (mul_34_17_n_11600 | mul_34_17_n_2025));
 assign mul_34_17_n_3928 = ((mul_34_17_n_1744 | mul_34_17_n_2360) & (mul_34_17_n_11600 | mul_34_17_n_1872));
 assign mul_34_17_n_3927 = (mul_34_17_n_2940 ^ mul_34_17_n_2829);
 assign mul_34_17_n_3926 = ~((mul_34_17_n_681 & mul_34_17_n_852) | (mul_34_17_n_2928 & mul_34_17_n_848));
 assign mul_34_17_n_3925 = ((mul_34_17_n_672 | mul_34_17_n_1050) & (mul_34_17_n_11552 | mul_34_17_n_1026));
 assign mul_34_17_n_3924 = ~((mul_34_17_n_1755 & mul_34_17_n_2431) | (mul_34_17_n_2898 & mul_34_17_n_2385));
 assign mul_34_17_n_3923 = ((mul_34_17_n_664 | mul_34_17_n_1270) & (mul_34_17_n_11564 | mul_34_17_n_1282));
 assign mul_34_17_n_3922 = ((mul_34_17_n_1755 & mul_34_17_n_2145) | (mul_34_17_n_2898 & mul_34_17_n_2088));
 assign mul_34_17_n_3920 = ((mul_34_17_n_673 & mul_34_17_n_1062) | (mul_34_17_n_2920 & mul_34_17_n_1044));
 assign mul_34_17_n_3919 = ((mul_34_17_n_663 & mul_34_17_n_1308) | (mul_34_17_n_2910 & mul_34_17_n_1330));
 assign mul_34_17_n_3917 = ((mul_34_17_n_1750 | mul_34_17_n_2583) & (mul_34_17_n_11612 | mul_34_17_n_2678));
 assign mul_34_17_n_3916 = ((mul_34_17_n_672 | mul_34_17_n_1030) & (mul_34_17_n_11552 | mul_34_17_n_1050));
 assign mul_34_17_n_3915 = ((mul_34_17_n_656 | mul_34_17_n_1531) & (mul_34_17_n_11576 | mul_34_17_n_1565));
 assign mul_34_17_n_3914 = ~((mul_34_17_n_674 | mul_34_17_n_1005) & (mul_34_17_n_11549 | mul_34_17_n_985));
 assign mul_34_17_n_3913 = ((mul_34_17_n_1740 | mul_34_17_n_2322) & (mul_34_17_n_11603 | mul_34_17_n_2057));
 assign mul_34_17_n_3912 = ((mul_34_17_n_1749 & mul_34_17_n_2569) | (mul_34_17_n_2890 & mul_34_17_n_2247));
 assign mul_34_17_n_3911 = ~((mul_34_17_n_663 & mul_34_17_n_1322) | (mul_34_17_n_2910 & mul_34_17_n_1338));
 assign mul_34_17_n_3910 = ~((mul_34_17_n_681 & mul_34_17_n_835) | (mul_34_17_n_2928 & mul_34_17_n_841));
 assign mul_34_17_n_3909 = ((mul_34_17_n_1754 | mul_34_17_n_2420) & (mul_34_17_n_11585 | mul_34_17_n_2296));
 assign mul_34_17_n_3908 = ~((mul_34_17_n_663 & mul_34_17_n_1325) | (mul_34_17_n_2910 & mul_34_17_n_1352));
 assign mul_34_17_n_3907 = ((mul_34_17_n_658 | mul_34_17_n_1468) & (mul_34_17_n_11573 | mul_34_17_n_1483));
 assign mul_34_17_n_3906 = ((mul_34_17_n_682 | mul_34_17_n_829) & (mul_34_17_n_11537 | mul_34_17_n_809));
 assign mul_34_17_n_3904 = ((mul_34_17_n_1752 | mul_34_17_n_2020) & (mul_34_17_n_11615 | mul_34_17_n_2242));
 assign mul_34_17_n_3903 = ((mul_34_17_n_668 | mul_34_17_n_1170) & (mul_34_17_n_11558 | mul_34_17_n_1142));
 assign mul_34_17_n_3902 = ((mul_34_17_n_1736 | mul_34_17_n_2215) & (mul_34_17_n_11591 | mul_34_17_n_1979));
 assign mul_34_17_n_3900 = ~((mul_34_17_n_682 | mul_34_17_n_809) & (mul_34_17_n_11537 | mul_34_17_n_816));
 assign mul_34_17_n_3899 = ~((mul_34_17_n_667 & mul_34_17_n_1224) | (mul_34_17_n_2914 & mul_34_17_n_1210));
 assign mul_34_17_n_3898 = ((mul_34_17_n_680 | mul_34_17_n_844) & (mul_34_17_n_11540 | mul_34_17_n_862));
 assign mul_34_17_n_3896 = ((mul_34_17_n_656 | mul_34_17_n_1524) & (mul_34_17_n_11576 | mul_34_17_n_1534));
 assign mul_34_17_n_3895 = ((mul_34_17_n_680 | mul_34_17_n_845) & (mul_34_17_n_11540 | mul_34_17_n_850));
 assign mul_34_17_n_3894 = ((mul_34_17_n_688 | mul_34_17_n_725) & (mul_34_17_n_11528 | mul_34_17_n_842));
 assign mul_34_17_n_3893 = ((mul_34_17_n_684 | mul_34_17_n_793) & (mul_34_17_n_11534 | mul_34_17_n_774));
 assign mul_34_17_n_3892 = ((mul_34_17_n_1734 | mul_34_17_n_2633) & (mul_34_17_n_11588 | mul_34_17_n_2494));
 assign mul_34_17_n_3891 = ((mul_34_17_n_1738 | mul_34_17_n_2458) & (mul_34_17_n_11606 | mul_34_17_n_2263));
 assign mul_34_17_n_3889 = ((mul_34_17_n_674 | mul_34_17_n_974) & (mul_34_17_n_11549 | mul_34_17_n_978));
 assign mul_34_17_n_3888 = ((mul_34_17_n_1734 | mul_34_17_n_2441) & (mul_34_17_n_11588 | mul_34_17_n_2173));
 assign mul_34_17_n_3887 = ((mul_34_17_n_1734 | mul_34_17_n_2701) & (mul_34_17_n_11588 | mul_34_17_n_2264));
 assign mul_34_17_n_3886 = ((mul_34_17_n_1736 | mul_34_17_n_2208) & (mul_34_17_n_11591 | mul_34_17_n_2511));
 assign mul_34_17_n_3885 = ((mul_34_17_n_672 | mul_34_17_n_1048) & (mul_34_17_n_11552 | mul_34_17_n_1028));
 assign mul_34_17_n_3884 = ((mul_34_17_n_682 | mul_34_17_n_816) & (mul_34_17_n_11537 | mul_34_17_n_823));
 assign mul_34_17_n_3883 = ~((mul_34_17_n_664 | mul_34_17_n_1288) & (mul_34_17_n_11564 | mul_34_17_n_1284));
 assign mul_34_17_n_3882 = ((mul_34_17_n_672 | mul_34_17_n_1023) & (mul_34_17_n_11552 | mul_34_17_n_1056));
 assign mul_34_17_n_3881 = ~((mul_34_17_n_1743 & mul_34_17_n_2282) | (mul_34_17_n_2882 & mul_34_17_n_1863));
 assign mul_34_17_n_3880 = ~((mul_34_17_n_1755 & mul_34_17_n_1858) | (mul_34_17_n_2898 & mul_34_17_n_1882));
 assign mul_34_17_n_3879 = ~((mul_34_17_n_1746 | mul_34_17_n_2184) & (mul_34_17_n_11652 | mul_34_17_n_2367));
 assign mul_34_17_n_3878 = ((mul_34_17_n_676 | mul_34_17_n_958) & (mul_34_17_n_11546 | mul_34_17_n_927));
 assign mul_34_17_n_3877 = ((mul_34_17_n_664 | mul_34_17_n_1274) & (mul_34_17_n_11564 | mul_34_17_n_1293));
 assign mul_34_17_n_3876 = ((mul_34_17_n_1750 | mul_34_17_n_2675) & (mul_34_17_n_11612 | mul_34_17_n_2364));
 assign mul_34_17_n_3875 = ((mul_34_17_n_680 | mul_34_17_n_867) & (mul_34_17_n_11540 | mul_34_17_n_834));
 assign mul_34_17_n_3874 = ((mul_34_17_n_1738 | mul_34_17_n_1856) & (mul_34_17_n_11606 | mul_34_17_n_2188));
 assign mul_34_17_n_3873 = ((mul_34_17_n_1752 | mul_34_17_n_2199) & (mul_34_17_n_11615 | mul_34_17_n_1929));
 assign mul_34_17_n_3872 = ~((mul_34_17_n_1753 & mul_34_17_n_2259) | (mul_34_17_n_2878 & mul_34_17_n_2444));
 assign mul_34_17_n_3871 = ((mul_34_17_n_660 | mul_34_17_n_1416) & (mul_34_17_n_11570 | mul_34_17_n_1398));
 assign mul_34_17_n_3870 = ((mul_34_17_n_666 | mul_34_17_n_1208) & (mul_34_17_n_11561 | mul_34_17_n_1201));
 assign mul_34_17_n_3869 = ((mul_34_17_n_668 | mul_34_17_n_1168) & (mul_34_17_n_11558 | mul_34_17_n_1164));
 assign mul_34_17_n_3868 = ((mul_34_17_n_1737 & mul_34_17_n_2411) | (mul_34_17_n_2894 & mul_34_17_n_1962));
 assign mul_34_17_n_3867 = ~((mul_34_17_n_1755 & mul_34_17_n_2396) | (mul_34_17_n_2898 & mul_34_17_n_2145));
 assign mul_34_17_n_3866 = ((mul_34_17_n_1754 | mul_34_17_n_2608) & (mul_34_17_n_11585 | mul_34_17_n_2445));
 assign mul_34_17_n_3865 = ((mul_34_17_n_1750 | mul_34_17_n_2220) & (mul_34_17_n_11612 | mul_34_17_n_2437));
 assign mul_34_17_n_3864 = ((mul_34_17_n_670 | mul_34_17_n_1074) & (mul_34_17_n_11555 | mul_34_17_n_1103));
 assign mul_34_17_n_3862 = ((mul_34_17_n_1756 | mul_34_17_n_866) & (mul_34_17_n_11582 | mul_34_17_n_1176));
 assign mul_34_17_n_3861 = ~((mul_34_17_n_664 | mul_34_17_n_1255) & (mul_34_17_n_11564 | mul_34_17_n_1273));
 assign mul_34_17_n_3859 = ((mul_34_17_n_660 | mul_34_17_n_1430) & (mul_34_17_n_11570 | mul_34_17_n_1393));
 assign mul_34_17_n_3858 = ((mul_34_17_n_1744 | mul_34_17_n_2164) & (mul_34_17_n_11600 | mul_34_17_n_2529));
 assign mul_34_17_n_3042 = ~(mul_34_17_n_2993 | mul_34_17_n_2744);
 assign mul_34_17_n_3856 = ((mul_34_17_n_1750 | mul_34_17_n_2085) & (mul_34_17_n_11612 | mul_34_17_n_2606));
 assign mul_34_17_n_3855 = ((mul_34_17_n_1756 | mul_34_17_n_1677) & (mul_34_17_n_11582 | mul_34_17_n_1758));
 assign mul_34_17_n_3854 = ~((mul_34_17_n_1743 & mul_34_17_n_2275) | (mul_34_17_n_2882 & mul_34_17_n_2118));
 assign mul_34_17_n_3853 = ~((mul_34_17_n_1747 & mul_34_17_n_2562) | (mul_34_17_n_11593 & mul_34_17_n_2028));
 assign mul_34_17_n_3852 = ~((mul_34_17_n_1754 | mul_34_17_n_1906) & (mul_34_17_n_11585 | mul_34_17_n_2154));
 assign mul_34_17_n_3850 = ~((mul_34_17_n_678 | mul_34_17_n_899) & (mul_34_17_n_11543 | mul_34_17_n_878));
 assign mul_34_17_n_3848 = ~((mul_34_17_n_1744 | mul_34_17_n_2034) & (mul_34_17_n_11600 | mul_34_17_n_2329));
 assign mul_34_17_n_3847 = ~((mul_34_17_n_1745 & mul_34_17_n_2689) | (mul_34_17_n_2888 & mul_34_17_n_2258));
 assign mul_34_17_n_3845 = ((mul_34_17_n_684 | mul_34_17_n_778) & (mul_34_17_n_11534 | mul_34_17_n_793));
 assign mul_34_17_n_3844 = ~((mul_34_17_n_663 & mul_34_17_n_1360) | (mul_34_17_n_2910 & mul_34_17_n_1372));
 assign mul_34_17_n_3843 = ((mul_34_17_n_1736 | mul_34_17_n_2394) & (mul_34_17_n_11591 | mul_34_17_n_2347));
 assign mul_34_17_n_3842 = ~((mul_34_17_n_1739 & mul_34_17_n_2123) | (mul_34_17_n_2884 & mul_34_17_n_2639));
 assign mul_34_17_n_3841 = ((mul_34_17_n_676 | mul_34_17_n_931) & (mul_34_17_n_11546 | mul_34_17_n_929));
 assign mul_34_17_n_3840 = ((mul_34_17_n_688 | mul_34_17_n_726) & (mul_34_17_n_11528 | mul_34_17_n_1702));
 assign mul_34_17_n_3839 = ((mul_34_17_n_1752 | mul_34_17_n_2042) & (mul_34_17_n_11615 | mul_34_17_n_2262));
 assign mul_34_17_n_3837 = ~((mul_34_17_n_1747 & mul_34_17_n_2472) | (mul_34_17_n_11593 & mul_34_17_n_1945));
 assign mul_34_17_n_3836 = ((mul_34_17_n_678 | mul_34_17_n_904) & (mul_34_17_n_11543 | mul_34_17_n_887));
 assign mul_34_17_n_3835 = ~((mul_34_17_n_1753 & mul_34_17_n_2680) | (mul_34_17_n_2878 & mul_34_17_n_1840));
 assign mul_34_17_n_3834 = ((mul_34_17_n_1735 & mul_34_17_n_1926) | (mul_34_17_n_2896 & mul_34_17_n_2062));
 assign mul_34_17_n_3833 = ~((mul_34_17_n_1745 & mul_34_17_n_2104) | (mul_34_17_n_2888 & mul_34_17_n_2686));
 assign mul_34_17_n_3832 = ((mul_34_17_n_1752 | mul_34_17_n_2650) & (mul_34_17_n_11615 | mul_34_17_n_2400));
 assign mul_34_17_n_3831 = ((mul_34_17_n_1748 | mul_34_17_n_2121) & (mul_34_17_n_11597 | mul_34_17_n_1869));
 assign mul_34_17_n_3830 = ((mul_34_17_n_1744 | mul_34_17_n_2267) & (mul_34_17_n_11600 | mul_34_17_n_2403));
 assign mul_34_17_n_3829 = ((mul_34_17_n_1756 | mul_34_17_n_1681) & (mul_34_17_n_11582 | mul_34_17_n_1576));
 assign mul_34_17_n_3828 = ((mul_34_17_n_1737 & mul_34_17_n_2221) | (mul_34_17_n_2894 & mul_34_17_n_2573));
 assign mul_34_17_n_3827 = ((mul_34_17_n_682 | mul_34_17_n_810) & (mul_34_17_n_11537 | mul_34_17_n_808));
 assign mul_34_17_n_3826 = ((mul_34_17_n_686 | mul_34_17_n_1112) & (mul_34_17_n_11531 | mul_34_17_n_735));
 assign mul_34_17_n_3825 = ~((mul_34_17_n_668 | mul_34_17_n_1140) & (mul_34_17_n_11558 | mul_34_17_n_1182));
 assign mul_34_17_n_3824 = ((mul_34_17_n_1746 | mul_34_17_n_1946) & (mul_34_17_n_11683 | mul_34_17_n_2147));
 assign mul_34_17_n_3822 = ((mul_34_17_n_1746 | mul_34_17_n_2283) & (mul_34_17_n_11685 | mul_34_17_n_2519));
 assign mul_34_17_n_3821 = ((mul_34_17_n_664 | mul_34_17_n_1256) & (mul_34_17_n_11564 | mul_34_17_n_1254));
 assign mul_34_17_n_3819 = ((mul_34_17_n_678 | mul_34_17_n_896) & (mul_34_17_n_11543 | mul_34_17_n_879));
 assign mul_34_17_n_3818 = ~((mul_34_17_n_1757 & mul_34_17_n_1671) | (mul_34_17_n_2900 & mul_34_17_n_1683));
 assign mul_34_17_n_3817 = ((mul_34_17_n_658 | mul_34_17_n_1471) & (mul_34_17_n_11573 | mul_34_17_n_1451));
 assign mul_34_17_n_3816 = ((mul_34_17_n_662 | mul_34_17_n_1313) & (mul_34_17_n_11567 | mul_34_17_n_1373));
 assign mul_34_17_n_3815 = ((mul_34_17_n_1742 | mul_34_17_n_2160) & (mul_34_17_n_11609 | mul_34_17_n_2166));
 assign mul_34_17_n_3814 = ((mul_34_17_n_1736 | mul_34_17_n_2525) & (mul_34_17_n_11591 | mul_34_17_n_2066));
 assign mul_34_17_n_3813 = ((mul_34_17_n_678 | mul_34_17_n_887) & (mul_34_17_n_11543 | mul_34_17_n_899));
 assign mul_34_17_n_3812 = ((mul_34_17_n_680 | mul_34_17_n_851) & (mul_34_17_n_11540 | mul_34_17_n_872));
 assign mul_34_17_n_3811 = ((mul_34_17_n_676 | mul_34_17_n_920) & (mul_34_17_n_11546 | mul_34_17_n_950));
 assign mul_34_17_n_3810 = ((mul_34_17_n_1742 | mul_34_17_n_2425) & (mul_34_17_n_11609 | mul_34_17_n_2058));
 assign mul_34_17_n_3809 = ~((mul_34_17_n_657 & mul_34_17_n_1580) | (mul_34_17_n_2904 & mul_34_17_n_1535));
 assign mul_34_17_n_3808 = ~((mul_34_17_n_655 & mul_34_17_n_1654) | (mul_34_17_n_2902 & mul_34_17_n_1661));
 assign mul_34_17_n_3807 = ~((mul_34_17_n_1734 | mul_34_17_n_2060) & (mul_34_17_n_11588 | mul_34_17_n_2368));
 assign mul_34_17_n_3806 = ~((mul_34_17_n_1749 & mul_34_17_n_2235) | (mul_34_17_n_2890 & mul_34_17_n_2011));
 assign mul_34_17_n_3804 = ((mul_34_17_n_666 | mul_34_17_n_1192) & (mul_34_17_n_11561 | mul_34_17_n_1198));
 assign mul_34_17_n_3802 = ((mul_34_17_n_1754 | mul_34_17_n_2055) & (mul_34_17_n_11585 | mul_34_17_n_1921));
 assign mul_34_17_n_3801 = ~((mul_34_17_n_665 & mul_34_17_n_1287) | (mul_34_17_n_2912 & mul_34_17_n_1259));
 assign mul_34_17_n_3800 = ((mul_34_17_n_1738 | mul_34_17_n_2053) & (mul_34_17_n_11606 | mul_34_17_n_2052));
 assign mul_34_17_n_3799 = ~((mul_34_17_n_673 & mul_34_17_n_1039) | (mul_34_17_n_2920 & mul_34_17_n_1022));
 assign mul_34_17_n_3798 = ((mul_34_17_n_668 | mul_34_17_n_1182) & (mul_34_17_n_11558 | mul_34_17_n_1133));
 assign mul_34_17_n_3797 = ~((mul_34_17_n_659 & mul_34_17_n_1497) | (mul_34_17_n_2906 & mul_34_17_n_1464));
 assign mul_34_17_n_3796 = ((mul_34_17_n_1734 | mul_34_17_n_2688) & (mul_34_17_n_11588 | mul_34_17_n_2683));
 assign mul_34_17_n_3795 = ~((mul_34_17_n_677 & mul_34_17_n_940) | (mul_34_17_n_2924 & mul_34_17_n_967));
 assign mul_34_17_n_3794 = ~((mul_34_17_n_669 & mul_34_17_n_1184) | (mul_34_17_n_2916 & mul_34_17_n_1139));
 assign mul_34_17_n_3793 = ((mul_34_17_n_1756 | mul_34_17_n_1762) & (mul_34_17_n_11582 | mul_34_17_n_1775));
 assign mul_34_17_n_3792 = ~((mul_34_17_n_1745 & mul_34_17_n_2391) | (mul_34_17_n_2888 & mul_34_17_n_2205));
 assign mul_34_17_n_3791 = ((mul_34_17_n_666 | mul_34_17_n_1191) & (mul_34_17_n_11561 | mul_34_17_n_1225));
 assign mul_34_17_n_3790 = ~((mul_34_17_n_1745 & mul_34_17_n_2177) | (mul_34_17_n_2888 & mul_34_17_n_2597));
 assign mul_34_17_n_3789 = ~((mul_34_17_n_667 & mul_34_17_n_1246) | (mul_34_17_n_2914 & mul_34_17_n_1228));
 assign mul_34_17_n_3788 = ~((mul_34_17_n_1751 & mul_34_17_n_2036) | (mul_34_17_n_2880 & mul_34_17_n_2033));
 assign mul_34_17_n_3787 = ((mul_34_17_n_1752 | mul_34_17_n_2172) & (mul_34_17_n_11615 | mul_34_17_n_2068));
 assign mul_34_17_n_3786 = ~((mul_34_17_n_1743 & mul_34_17_n_2240) | (mul_34_17_n_2882 & mul_34_17_n_2249));
 assign mul_34_17_n_3785 = ((mul_34_17_n_1748 | mul_34_17_n_2549) & (mul_34_17_n_11597 | mul_34_17_n_2006));
 assign mul_34_17_n_3784 = ~((mul_34_17_n_668 | mul_34_17_n_1133) & (mul_34_17_n_11558 | mul_34_17_n_1143));
 assign mul_34_17_n_3783 = ((mul_34_17_n_1734 | mul_34_17_n_2416) & (mul_34_17_n_11588 | mul_34_17_n_2060));
 assign mul_34_17_n_3782 = ((mul_34_17_n_1752 | mul_34_17_n_2022) & (mul_34_17_n_11615 | mul_34_17_n_2469));
 assign mul_34_17_n_3781 = ((mul_34_17_n_674 | mul_34_17_n_984) & (mul_34_17_n_11549 | mul_34_17_n_971));
 assign mul_34_17_n_3779 = ((mul_34_17_n_1754 | mul_34_17_n_1950) & (mul_34_17_n_11585 | mul_34_17_n_2055));
 assign mul_34_17_n_3778 = ~((mul_34_17_n_658 | mul_34_17_n_1465) & (mul_34_17_n_11573 | mul_34_17_n_1505));
 assign mul_34_17_n_3776 = ((mul_34_17_n_1740 | mul_34_17_n_2099) & (mul_34_17_n_11603 | mul_34_17_n_2336));
 assign mul_34_17_n_3775 = ~((mul_34_17_n_1752 | mul_34_17_n_2012) & (mul_34_17_n_11615 | mul_34_17_n_2307));
 assign mul_34_17_n_3774 = ~((mul_34_17_n_1745 & mul_34_17_n_2274) | (mul_34_17_n_2888 & mul_34_17_n_2382));
 assign mul_34_17_n_3772 = ((mul_34_17_n_1736 | mul_34_17_n_2380) & (mul_34_17_n_11591 | mul_34_17_n_2551));
 assign mul_34_17_n_3771 = ((mul_34_17_n_1744 | mul_34_17_n_2017) & (mul_34_17_n_11600 | mul_34_17_n_2693));
 assign mul_34_17_n_3770 = ~((mul_34_17_n_672 | mul_34_17_n_1021) & (mul_34_17_n_11552 | mul_34_17_n_1052));
 assign mul_34_17_n_3769 = ((mul_34_17_n_1749 & mul_34_17_n_2044) | (mul_34_17_n_2890 & mul_34_17_n_2665));
 assign mul_34_17_n_3768 = ~((mul_34_17_n_667 & mul_34_17_n_1199) | (mul_34_17_n_2914 & mul_34_17_n_1247));
 assign mul_34_17_n_3766 = ((mul_34_17_n_1748 | mul_34_17_n_2076) & (mul_34_17_n_11597 | mul_34_17_n_1904));
 assign mul_34_17_n_3765 = ((mul_34_17_n_1747 & mul_34_17_n_2638) | (mul_34_17_n_11593 & mul_34_17_n_1886));
 assign mul_34_17_n_3764 = ((mul_34_17_n_668 | mul_34_17_n_1135) & (mul_34_17_n_11558 | mul_34_17_n_1129));
 assign mul_34_17_n_3762 = ((mul_34_17_n_668 | mul_34_17_n_1131) & (mul_34_17_n_11558 | mul_34_17_n_1183));
 assign mul_34_17_n_3761 = ((mul_34_17_n_682 | mul_34_17_n_817) & (mul_34_17_n_11537 | mul_34_17_n_801));
 assign mul_34_17_n_3760 = ~((mul_34_17_n_661 & mul_34_17_n_1413) | (mul_34_17_n_2908 & mul_34_17_n_1409));
 assign mul_34_17_n_3759 = ((mul_34_17_n_1750 | mul_34_17_n_2508) & (mul_34_17_n_11612 | mul_34_17_n_2603));
 assign mul_34_17_n_3758 = ((mul_34_17_n_656 | mul_34_17_n_1549) & (mul_34_17_n_11576 | mul_34_17_n_1566));
 assign mul_34_17_n_3757 = ((mul_34_17_n_676 | mul_34_17_n_953) & (mul_34_17_n_11546 | mul_34_17_n_926));
 assign mul_34_17_n_3756 = ((mul_34_17_n_1753 & mul_34_17_n_2594) | (mul_34_17_n_2878 & mul_34_17_n_2217));
 assign mul_34_17_n_3755 = ((mul_34_17_n_1752 | mul_34_17_n_1969) & (mul_34_17_n_11615 | mul_34_17_n_1944));
 assign mul_34_17_n_3754 = ~((mul_34_17_n_657 & mul_34_17_n_1525) | (mul_34_17_n_2904 & mul_34_17_n_1582));
 assign mul_34_17_n_3753 = ((mul_34_17_n_658 | mul_34_17_n_1463) & (mul_34_17_n_11573 | mul_34_17_n_1467));
 assign mul_34_17_n_3752 = ~((mul_34_17_n_663 & mul_34_17_n_1329) | (mul_34_17_n_2910 & mul_34_17_n_1312));
 assign mul_34_17_n_3751 = ((mul_34_17_n_1748 | mul_34_17_n_1898) & (mul_34_17_n_11597 | mul_34_17_n_2111));
 assign mul_34_17_n_3750 = ((mul_34_17_n_1742 | mul_34_17_n_2348) & (mul_34_17_n_11609 | mul_34_17_n_1988));
 assign mul_34_17_n_3749 = ((mul_34_17_n_655 & mul_34_17_n_1660) | (mul_34_17_n_2902 & mul_34_17_n_1597));
 assign mul_34_17_n_3748 = ((mul_34_17_n_658 | mul_34_17_n_1467) & (mul_34_17_n_11573 | mul_34_17_n_1500));
 assign mul_34_17_n_3747 = ((mul_34_17_n_662 | mul_34_17_n_1348) & (mul_34_17_n_11567 | mul_34_17_n_1316));
 assign mul_34_17_n_3746 = ((mul_34_17_n_1742 | mul_34_17_n_1961) & (mul_34_17_n_11609 | mul_34_17_n_2183));
 assign mul_34_17_n_3744 = ((mul_34_17_n_660 | mul_34_17_n_1401) & (mul_34_17_n_11570 | mul_34_17_n_1381));
 assign mul_34_17_n_3743 = ~((mul_34_17_n_1743 & mul_34_17_n_2321) | (mul_34_17_n_2882 & mul_34_17_n_1956));
 assign mul_34_17_n_3742 = ((mul_34_17_n_1750 | mul_34_17_n_1954) & (mul_34_17_n_11612 | mul_34_17_n_2448));
 assign mul_34_17_n_3741 = ((mul_34_17_n_678 | mul_34_17_n_891) & (mul_34_17_n_11543 | mul_34_17_n_908));
 assign mul_34_17_n_3740 = ((mul_34_17_n_670 | mul_34_17_n_1100) & (mul_34_17_n_11555 | mul_34_17_n_1084));
 assign mul_34_17_n_3739 = ((mul_34_17_n_1742 | mul_34_17_n_2191) & (mul_34_17_n_11609 | mul_34_17_n_2471));
 assign mul_34_17_n_3738 = ~((mul_34_17_n_659 & mul_34_17_n_1477) | (mul_34_17_n_2906 & mul_34_17_n_1480));
 assign mul_34_17_n_3737 = ((mul_34_17_n_664 | mul_34_17_n_1252) & (mul_34_17_n_11564 | mul_34_17_n_1275));
 assign mul_34_17_n_3736 = ~((mul_34_17_n_1745 & mul_34_17_n_2682) | (mul_34_17_n_2888 & mul_34_17_n_2115));
 assign mul_34_17_n_3735 = ((mul_34_17_n_675 & mul_34_17_n_998) | (mul_34_17_n_2922 & mul_34_17_n_991));
 assign mul_34_17_n_3734 = ((mul_34_17_n_1740 | mul_34_17_n_2438) & (mul_34_17_n_11603 | mul_34_17_n_2231));
 assign mul_34_17_n_3733 = ((mul_34_17_n_1754 | mul_34_17_n_2296) & (mul_34_17_n_11585 | mul_34_17_n_1967));
 assign mul_34_17_n_3732 = ~((mul_34_17_n_1743 & mul_34_17_n_2334) | (mul_34_17_n_2882 & mul_34_17_n_2609));
 assign mul_34_17_n_3731 = ((mul_34_17_n_662 | mul_34_17_n_1356) & (mul_34_17_n_11567 | mul_34_17_n_1365));
 assign mul_34_17_n_3730 = ((mul_34_17_n_1738 | mul_34_17_n_1696) & (mul_34_17_n_11606 | mul_34_17_n_2504));
 assign mul_34_17_n_3729 = ((mul_34_17_n_682 | mul_34_17_n_820) & (mul_34_17_n_11537 | mul_34_17_n_826));
 assign mul_34_17_n_3728 = ~((mul_34_17_n_1735 & mul_34_17_n_1942) | (mul_34_17_n_2896 & mul_34_17_n_2131));
 assign mul_34_17_n_3727 = ((mul_34_17_n_1742 | mul_34_17_n_2479) & (mul_34_17_n_11609 | mul_34_17_n_2191));
 assign mul_34_17_n_3726 = ((mul_34_17_n_1742 | mul_34_17_n_2229) & (mul_34_17_n_11609 | mul_34_17_n_2265));
 assign mul_34_17_n_3725 = ((mul_34_17_n_1746 | mul_34_17_n_2439) & (mul_34_17_n_11649 | mul_34_17_n_2297));
 assign mul_34_17_n_3724 = ((mul_34_17_n_654 | mul_34_17_n_1638) & (mul_34_17_n_11579 | mul_34_17_n_1591));
 assign mul_34_17_n_3723 = ~((mul_34_17_n_665 & mul_34_17_n_1297) | (mul_34_17_n_2912 & mul_34_17_n_1265));
 assign mul_34_17_n_3721 = ((mul_34_17_n_1740 | mul_34_17_n_2514) & (mul_34_17_n_11603 | mul_34_17_n_2405));
 assign mul_34_17_n_3720 = ((mul_34_17_n_1750 | mul_34_17_n_2500) & (mul_34_17_n_11612 | mul_34_17_n_2065));
 assign mul_34_17_n_3719 = ~((mul_34_17_n_677 & mul_34_17_n_942) | (mul_34_17_n_2924 & mul_34_17_n_928));
 assign mul_34_17_n_3718 = ((mul_34_17_n_1750 | mul_34_17_n_1963) & (mul_34_17_n_11612 | mul_34_17_n_2330));
 assign mul_34_17_n_3717 = ((mul_34_17_n_656 | mul_34_17_n_1527) & (mul_34_17_n_11576 | mul_34_17_n_1575));
 assign mul_34_17_n_3716 = ((mul_34_17_n_1746 | mul_34_17_n_2147) & (mul_34_17_n_11663 | mul_34_17_n_2313));
 assign mul_34_17_n_3715 = ~((mul_34_17_n_1738 | mul_34_17_n_1911) & (mul_34_17_n_11606 | mul_34_17_n_1910));
 assign mul_34_17_n_3714 = ((mul_34_17_n_1742 | mul_34_17_n_2566) & (mul_34_17_n_11609 | mul_34_17_n_2462));
 assign mul_34_17_n_3713 = ((mul_34_17_n_1748 | mul_34_17_n_2029) & (mul_34_17_n_11597 | mul_34_17_n_2292));
 assign mul_34_17_n_3712 = ((mul_34_17_n_1740 | mul_34_17_n_2048) & (mul_34_17_n_11603 | mul_34_17_n_1985));
 assign mul_34_17_n_3711 = ((mul_34_17_n_658 | mul_34_17_n_1450) & (mul_34_17_n_11573 | mul_34_17_n_1508));
 assign mul_34_17_n_3710 = ~((mul_34_17_n_1752 | mul_34_17_n_2605) & (mul_34_17_n_11615 | mul_34_17_n_1915));
 assign mul_34_17_n_3709 = ((mul_34_17_n_1754 | mul_34_17_n_2610) & (mul_34_17_n_11585 | mul_34_17_n_1937));
 assign mul_34_17_n_3708 = ((mul_34_17_n_1752 | mul_34_17_n_2677) & (mul_34_17_n_11615 | mul_34_17_n_1874));
 assign mul_34_17_n_3707 = ((mul_34_17_n_1734 | mul_34_17_n_1909) & (mul_34_17_n_11588 | mul_34_17_n_2167));
 assign mul_34_17_n_3706 = ((mul_34_17_n_1736 | mul_34_17_n_2674) & (mul_34_17_n_11591 | mul_34_17_n_1932));
 assign mul_34_17_n_3705 = ((mul_34_17_n_660 | mul_34_17_n_1387) & (mul_34_17_n_11570 | mul_34_17_n_1375));
 assign mul_34_17_n_3704 = ((mul_34_17_n_1736 | mul_34_17_n_1891) & (mul_34_17_n_11591 | mul_34_17_n_2550));
 assign mul_34_17_n_3703 = ~((mul_34_17_n_679 & mul_34_17_n_913) | (mul_34_17_n_2926 & mul_34_17_n_889));
 assign mul_34_17_n_3701 = ((mul_34_17_n_664 | mul_34_17_n_1267) & (mul_34_17_n_11564 | mul_34_17_n_1252));
 assign mul_34_17_n_3700 = ((mul_34_17_n_658 | mul_34_17_n_1505) & (mul_34_17_n_11573 | mul_34_17_n_1496));
 assign mul_34_17_n_3699 = ((mul_34_17_n_1752 | mul_34_17_n_2156) & (mul_34_17_n_11615 | mul_34_17_n_2605));
 assign mul_34_17_n_3698 = ((mul_34_17_n_1744 | mul_34_17_n_1872) & (mul_34_17_n_11600 | mul_34_17_n_2015));
 assign mul_34_17_n_3696 = ((mul_34_17_n_1748 | mul_34_17_n_1883) & (mul_34_17_n_11597 | mul_34_17_n_2538));
 assign mul_34_17_n_3694 = ((mul_34_17_n_1746 | mul_34_17_n_2189) & (mul_34_17_n_11644 | mul_34_17_n_2356));
 assign mul_34_17_n_3693 = ~((mul_34_17_n_1757 & mul_34_17_n_1003) | (mul_34_17_n_2900 & mul_34_17_n_1761));
 assign mul_34_17_n_3692 = ~((mul_34_17_n_1747 & mul_34_17_n_1878) | (mul_34_17_n_11593 & mul_34_17_n_2212));
 assign mul_34_17_n_3691 = ((mul_34_17_n_1755 & mul_34_17_n_2670) | (mul_34_17_n_2898 & mul_34_17_n_2219));
 assign mul_34_17_n_3690 = ~((mul_34_17_n_1736 | mul_34_17_n_2465) & (mul_34_17_n_11591 | mul_34_17_n_1891));
 assign mul_34_17_n_3689 = ((mul_34_17_n_1740 | mul_34_17_n_2079) & (mul_34_17_n_11603 | mul_34_17_n_2438));
 assign mul_34_17_n_3687 = ((mul_34_17_n_666 | mul_34_17_n_1232) & (mul_34_17_n_11561 | mul_34_17_n_1235));
 assign mul_34_17_n_3685 = ((mul_34_17_n_666 | mul_34_17_n_1221) & (mul_34_17_n_11561 | mul_34_17_n_1207));
 assign mul_34_17_n_3684 = ((mul_34_17_n_672 | mul_34_17_n_1052) & (mul_34_17_n_11552 | mul_34_17_n_1017));
 assign mul_34_17_n_3682 = ((mul_34_17_n_1752 | mul_34_17_n_1874) & (mul_34_17_n_11615 | mul_34_17_n_2156));
 assign mul_34_17_n_3681 = ~((mul_34_17_n_671 & mul_34_17_n_1091) | (mul_34_17_n_2918 & mul_34_17_n_1119));
 assign mul_34_17_n_3679 = ((mul_34_17_n_668 | mul_34_17_n_1143) & (mul_34_17_n_11558 | mul_34_17_n_1150));
 assign mul_34_17_n_3678 = ((mul_34_17_n_657 & mul_34_17_n_1585) | (mul_34_17_n_2904 & mul_34_17_n_1528));
 assign mul_34_17_n_3677 = ((mul_34_17_n_666 | mul_34_17_n_1229) & (mul_34_17_n_11561 | mul_34_17_n_1232));
 assign mul_34_17_n_3676 = ((mul_34_17_n_1750 | mul_34_17_n_2555) & (mul_34_17_n_11612 | mul_34_17_n_1857));
 assign mul_34_17_n_3675 = ((mul_34_17_n_674 | mul_34_17_n_987) & (mul_34_17_n_11549 | mul_34_17_n_999));
 assign mul_34_17_n_3674 = ((mul_34_17_n_654 | mul_34_17_n_1614) & (mul_34_17_n_11579 | mul_34_17_n_1594));
 assign mul_34_17_n_3673 = ((mul_34_17_n_678 | mul_34_17_n_895) & (mul_34_17_n_11543 | mul_34_17_n_914));
 assign mul_34_17_n_3672 = ~((mul_34_17_n_655 & mul_34_17_n_1604) | (mul_34_17_n_2902 & mul_34_17_n_1619));
 assign mul_34_17_n_3671 = ~((mul_34_17_n_1753 & mul_34_17_n_2217) | (mul_34_17_n_2878 & mul_34_17_n_2567));
 assign mul_34_17_n_3669 = ~((mul_34_17_n_1739 & mul_34_17_n_1971) | (mul_34_17_n_2884 & mul_34_17_n_2203));
 assign mul_34_17_n_3668 = ((mul_34_17_n_1749 & mul_34_17_n_2268) | (mul_34_17_n_2890 & mul_34_17_n_1850));
 assign mul_34_17_n_3667 = ((mul_34_17_n_1736 | mul_34_17_n_2293) & (mul_34_17_n_11591 | mul_34_17_n_1901));
 assign mul_34_17_n_3666 = ((mul_34_17_n_1735 & mul_34_17_n_2070) | (mul_34_17_n_2896 & mul_34_17_n_2082));
 assign mul_34_17_n_3665 = ((mul_34_17_n_656 | mul_34_17_n_1532) & (mul_34_17_n_11576 | mul_34_17_n_1587));
 assign mul_34_17_n_3664 = ((mul_34_17_n_688 | mul_34_17_n_706) & (mul_34_17_n_11528 | mul_34_17_n_703));
 assign mul_34_17_n_3662 = ((mul_34_17_n_656 | mul_34_17_n_1575) & (mul_34_17_n_11576 | mul_34_17_n_1563));
 assign mul_34_17_n_3661 = ((mul_34_17_n_664 | mul_34_17_n_1264) & (mul_34_17_n_11564 | mul_34_17_n_1271));
 assign mul_34_17_n_3660 = (mul_34_17_n_2739 ^ mul_34_17_n_2848);
 assign mul_34_17_n_3659 = ((mul_34_17_n_1734 | mul_34_17_n_2324) & (mul_34_17_n_11588 | mul_34_17_n_2646));
 assign mul_34_17_n_3658 = ((mul_34_17_n_674 | mul_34_17_n_1007) & (mul_34_17_n_11549 | mul_34_17_n_982));
 assign mul_34_17_n_3657 = ~((mul_34_17_n_1742 | mul_34_17_n_2462) & (mul_34_17_n_11609 | mul_34_17_n_2496));
 assign mul_34_17_n_3656 = ((mul_34_17_n_1746 | mul_34_17_n_2227) & (mul_34_17_n_11662 | mul_34_17_n_2320));
 assign mul_34_17_n_3655 = ((mul_34_17_n_1756 | mul_34_17_n_827) & (mul_34_17_n_11582 | mul_34_17_n_1342));
 assign mul_34_17_n_3654 = ((mul_34_17_n_1740 | mul_34_17_n_2139) & (mul_34_17_n_11603 | mul_34_17_n_2285));
 assign mul_34_17_n_3653 = ((mul_34_17_n_1736 | mul_34_17_n_2066) & (mul_34_17_n_11591 | mul_34_17_n_2536));
 assign mul_34_17_n_3652 = ((mul_34_17_n_658 | mul_34_17_n_1473) & (mul_34_17_n_11573 | mul_34_17_n_1468));
 assign mul_34_17_n_3651 = ((mul_34_17_n_658 | mul_34_17_n_1500) & (mul_34_17_n_11573 | mul_34_17_n_1450));
 assign mul_34_17_n_3650 = ((mul_34_17_n_1736 | mul_34_17_n_2511) & (mul_34_17_n_11591 | mul_34_17_n_2178));
 assign mul_34_17_n_3649 = ~((mul_34_17_n_1749 & mul_34_17_n_2291) | (mul_34_17_n_2890 & mul_34_17_n_2196));
 assign mul_34_17_n_3648 = ~((mul_34_17_n_1751 & mul_34_17_n_2581) | (mul_34_17_n_2880 & mul_34_17_n_2654));
 assign mul_34_17_n_3647 = ((mul_34_17_n_690 | mul_34_17_n_741) & (mul_34_17_n_11525 | mul_34_17_n_745));
 assign mul_34_17_n_3646 = ((mul_34_17_n_1746 | mul_34_17_n_2356) & (mul_34_17_n_11697 | mul_34_17_n_2168));
 assign mul_34_17_n_3645 = ((mul_34_17_n_1742 | mul_34_17_n_2155) & (mul_34_17_n_11609 | mul_34_17_n_2450));
 assign mul_34_17_n_3643 = ~((mul_34_17_n_677 & mul_34_17_n_932) | (mul_34_17_n_2924 & mul_34_17_n_923));
 assign mul_34_17_n_3642 = ((mul_34_17_n_654 | mul_34_17_n_1635) & (mul_34_17_n_11579 | mul_34_17_n_1616));
 assign mul_34_17_n_3641 = ~((mul_34_17_n_1755 & mul_34_17_n_2211) | (mul_34_17_n_2898 & mul_34_17_n_2077));
 assign mul_34_17_n_3640 = ~((mul_34_17_n_1753 & mul_34_17_n_2397) | (mul_34_17_n_2878 & mul_34_17_n_2146));
 assign mul_34_17_n_3639 = ~((mul_34_17_n_688 | mul_34_17_n_694) & (mul_34_17_n_11528 | mul_34_17_n_701));
 assign mul_34_17_n_3638 = ~((mul_34_17_n_655 & mul_34_17_n_1642) | (mul_34_17_n_2902 & mul_34_17_n_1634));
 assign mul_34_17_n_3637 = ((mul_34_17_n_1734 | mul_34_17_n_2061) & (mul_34_17_n_11588 | mul_34_17_n_2284));
 assign mul_34_17_n_3635 = ~((mul_34_17_n_1741 & mul_34_17_n_2094) | (mul_34_17_n_2886 & mul_34_17_n_2461));
 assign mul_34_17_n_3634 = ((mul_34_17_n_1747 & mul_34_17_n_2314) | (mul_34_17_n_11593 & mul_34_17_n_2423));
 assign mul_34_17_n_3633 = ((mul_34_17_n_686 | mul_34_17_n_735) & (mul_34_17_n_11531 | mul_34_17_n_704));
 assign mul_34_17_n_3632 = ((mul_34_17_n_688 | mul_34_17_n_700) & (mul_34_17_n_11528 | mul_34_17_n_723));
 assign mul_34_17_n_3630 = ~((mul_34_17_n_679 & mul_34_17_n_912) | (mul_34_17_n_2926 & mul_34_17_n_881));
 assign mul_34_17_n_3629 = ((mul_34_17_n_1738 | mul_34_17_n_2310) & (mul_34_17_n_11606 | mul_34_17_n_2595));
 assign mul_34_17_n_3628 = ~((mul_34_17_n_1737 & mul_34_17_n_2544) | (mul_34_17_n_2894 & mul_34_17_n_2393));
 assign mul_34_17_n_3626 = ~((mul_34_17_n_1747 & mul_34_17_n_2080) | (mul_34_17_n_11593 & mul_34_17_n_2404));
 assign mul_34_17_n_3625 = ((mul_34_17_n_668 | mul_34_17_n_1150) & (mul_34_17_n_11558 | mul_34_17_n_1168));
 assign mul_34_17_n_3624 = ~((mul_34_17_n_1739 & mul_34_17_n_2339) | (mul_34_17_n_2884 & mul_34_17_n_2572));
 assign mul_34_17_n_3623 = ~((mul_34_17_n_1739 & mul_34_17_n_2300) | (mul_34_17_n_2884 & mul_34_17_n_2130));
 assign mul_34_17_n_3622 = ~((mul_34_17_n_1741 & mul_34_17_n_1984) | (mul_34_17_n_2886 & mul_34_17_n_2616));
 assign mul_34_17_n_3621 = ~((mul_34_17_n_663 & mul_34_17_n_1332) | (mul_34_17_n_2910 & mul_34_17_n_1366));
 assign mul_34_17_n_3620 = ((mul_34_17_n_1748 | mul_34_17_n_2142) & (mul_34_17_n_11597 | mul_34_17_n_2533));
 assign mul_34_17_n_3619 = ((mul_34_17_n_1740 | mul_34_17_n_2236) & (mul_34_17_n_11603 | mul_34_17_n_2216));
 assign mul_34_17_n_3618 = ((mul_34_17_n_678 | mul_34_17_n_890) & (mul_34_17_n_11543 | mul_34_17_n_894));
 assign mul_34_17_n_3617 = ((mul_34_17_n_1740 | mul_34_17_n_2030) & (mul_34_17_n_11603 | mul_34_17_n_1859));
 assign mul_34_17_n_3616 = ((mul_34_17_n_662 | mul_34_17_n_1339) & (mul_34_17_n_11567 | mul_34_17_n_1353));
 assign mul_34_17_n_3614 = ((mul_34_17_n_668 | mul_34_17_n_1142) & (mul_34_17_n_11558 | mul_34_17_n_1171));
 assign mul_34_17_n_3612 = ((mul_34_17_n_1746 | mul_34_17_n_2241) & (mul_34_17_n_11693 | mul_34_17_n_2560));
 assign mul_34_17_n_3611 = ((mul_34_17_n_666 | mul_34_17_n_1231) & (mul_34_17_n_11561 | mul_34_17_n_1221));
 assign mul_34_17_n_3610 = ~((mul_34_17_n_673 & mul_34_17_n_1053) | (mul_34_17_n_2920 & mul_34_17_n_1031));
 assign mul_34_17_n_3609 = ((mul_34_17_n_682 | mul_34_17_n_824) & (mul_34_17_n_11537 | mul_34_17_n_820));
 assign mul_34_17_n_3608 = ((mul_34_17_n_658 | mul_34_17_n_1446) & (mul_34_17_n_11573 | mul_34_17_n_1449));
 assign mul_34_17_n_3607 = ((mul_34_17_n_1754 | mul_34_17_n_2232) & (mul_34_17_n_11585 | mul_34_17_n_2430));
 assign mul_34_17_n_3606 = ((mul_34_17_n_666 | mul_34_17_n_1217) & (mul_34_17_n_11561 | mul_34_17_n_1219));
 assign mul_34_17_n_3605 = ((mul_34_17_n_666 | mul_34_17_n_1205) & (mul_34_17_n_11561 | mul_34_17_n_1227));
 assign mul_34_17_n_3603 = ((mul_34_17_n_1748 | mul_34_17_n_1869) & (mul_34_17_n_11597 | mul_34_17_n_2492));
 assign mul_34_17_n_3602 = ((mul_34_17_n_1750 | mul_34_17_n_2456) & (mul_34_17_n_11612 | mul_34_17_n_1991));
 assign mul_34_17_n_3601 = ((mul_34_17_n_656 | mul_34_17_n_1542) & (mul_34_17_n_11576 | mul_34_17_n_1570));
 assign mul_34_17_n_3600 = ((mul_34_17_n_662 | mul_34_17_n_1326) & (mul_34_17_n_11567 | mul_34_17_n_1309));
 assign mul_34_17_n_3599 = ((mul_34_17_n_1746 | mul_34_17_n_2585) & (mul_34_17_n_11659 | mul_34_17_n_2663));
 assign mul_34_17_n_3598 = ((mul_34_17_n_688 | mul_34_17_n_752) & (mul_34_17_n_11528 | mul_34_17_n_1200));
 assign mul_34_17_n_3597 = ~((mul_34_17_n_1745 & mul_34_17_n_2545) | (mul_34_17_n_2888 & mul_34_17_n_2149));
 assign mul_34_17_n_3595 = ~((mul_34_17_n_1739 & mul_34_17_n_2395) | (mul_34_17_n_2884 & mul_34_17_n_2300));
 assign mul_34_17_n_3594 = ((mul_34_17_n_1752 | mul_34_17_n_2286) & (mul_34_17_n_11615 | mul_34_17_n_2199));
 assign mul_34_17_n_3592 = ~((mul_34_17_n_1743 & mul_34_17_n_2497) | (mul_34_17_n_2882 & mul_34_17_n_2301));
 assign mul_34_17_n_3590 = ((mul_34_17_n_654 | mul_34_17_n_1645) & (mul_34_17_n_11579 | mul_34_17_n_1655));
 assign mul_34_17_n_3588 = ~((mul_34_17_n_669 & mul_34_17_n_1152) | (mul_34_17_n_2916 & mul_34_17_n_1169));
 assign mul_34_17_n_3587 = ~((mul_34_17_n_1739 & mul_34_17_n_2354) | (mul_34_17_n_2884 & mul_34_17_n_1841));
 assign mul_34_17_n_3586 = ~((mul_34_17_n_661 & mul_34_17_n_1423) | (mul_34_17_n_2908 & mul_34_17_n_1415));
 assign mul_34_17_n_3585 = ~((mul_34_17_n_687 & mul_34_17_n_740) | (mul_34_17_n_2933 & mul_34_17_n_744));
 assign mul_34_17_n_3584 = ((mul_34_17_n_656 | mul_34_17_n_1522) & (mul_34_17_n_11576 | mul_34_17_n_1529));
 assign mul_34_17_n_3583 = ((mul_34_17_n_660 | mul_34_17_n_1392) & (mul_34_17_n_11570 | mul_34_17_n_1411));
 assign mul_34_17_n_3582 = ((mul_34_17_n_688 | mul_34_17_n_692) & (mul_34_17_n_11528 | mul_34_17_n_698));
 assign mul_34_17_n_3581 = ~((mul_34_17_n_670 | mul_34_17_n_1109) & (mul_34_17_n_11555 | mul_34_17_n_1071));
 assign mul_34_17_n_3580 = ~((mul_34_17_n_685 & mul_34_17_n_764) | (mul_34_17_n_2931 & mul_34_17_n_765));
 assign mul_34_17_n_3579 = ((mul_34_17_n_1737 & mul_34_17_n_2552) | (mul_34_17_n_2894 & mul_34_17_n_2631));
 assign mul_34_17_n_3578 = ((mul_34_17_n_1746 | mul_34_17_n_2152) & (mul_34_17_n_11686 | mul_34_17_n_2412));
 assign mul_34_17_n_3576 = ~((mul_34_17_n_1741 & mul_34_17_n_2331) | (mul_34_17_n_2886 & mul_34_17_n_2120));
 assign mul_34_17_n_3575 = ((mul_34_17_n_688 | mul_34_17_n_1266) & (mul_34_17_n_11528 | mul_34_17_n_752));
 assign mul_34_17_n_3574 = ((mul_34_17_n_1744 | mul_34_17_n_2421) & (mul_34_17_n_11600 | mul_34_17_n_2399));
 assign mul_34_17_n_3573 = ((mul_34_17_n_666 | mul_34_17_n_1238) & (mul_34_17_n_11561 | mul_34_17_n_1226));
 assign mul_34_17_n_3572 = ((mul_34_17_n_1740 | mul_34_17_n_2285) & (mul_34_17_n_11603 | mul_34_17_n_2099));
 assign mul_34_17_n_3571 = ((mul_34_17_n_1746 | mul_34_17_n_1864) & (mul_34_17_n_11696 | mul_34_17_n_2241));
 assign mul_34_17_n_3570 = ~((mul_34_17_n_669 & mul_34_17_n_1130) | (mul_34_17_n_2916 & mul_34_17_n_1141));
 assign mul_34_17_n_3568 = ~((mul_34_17_n_669 & mul_34_17_n_1132) | (mul_34_17_n_2916 & mul_34_17_n_1145));
 assign mul_34_17_n_3567 = ((mul_34_17_n_670 | mul_34_17_n_1088) & (mul_34_17_n_11555 | mul_34_17_n_1068));
 assign mul_34_17_n_3566 = ((mul_34_17_n_1750 | mul_34_17_n_2606) & (mul_34_17_n_11612 | mul_34_17_n_2387));
 assign mul_34_17_n_3565 = ~((mul_34_17_n_675 & mul_34_17_n_991) | (mul_34_17_n_2922 & mul_34_17_n_976));
 assign mul_34_17_n_3564 = ((mul_34_17_n_665 & mul_34_17_n_1294) | (mul_34_17_n_2912 & mul_34_17_n_1263));
 assign mul_34_17_n_3563 = ((mul_34_17_n_688 | mul_34_17_n_769) & (mul_34_17_n_11528 | mul_34_17_n_755));
 assign mul_34_17_n_3562 = ((mul_34_17_n_666 | mul_34_17_n_1236) & (mul_34_17_n_11561 | mul_34_17_n_1231));
 assign mul_34_17_n_3561 = ((mul_34_17_n_1747 & mul_34_17_n_2100) | (mul_34_17_n_11593 & mul_34_17_n_1865));
 assign mul_34_17_n_3560 = ((mul_34_17_n_666 | mul_34_17_n_1234) & (mul_34_17_n_11561 | mul_34_17_n_1203));
 assign mul_34_17_n_3559 = ~((mul_34_17_n_671 & mul_34_17_n_1083) | (mul_34_17_n_2918 & mul_34_17_n_1075));
 assign mul_34_17_n_3558 = ~((mul_34_17_n_1743 & mul_34_17_n_2695) | (mul_34_17_n_2882 & mul_34_17_n_2535));
 assign mul_34_17_n_3556 = ((mul_34_17_n_662 | mul_34_17_n_1321) & (mul_34_17_n_11567 | mul_34_17_n_1345));
 assign mul_34_17_n_3554 = ((mul_34_17_n_1742 | mul_34_17_n_2471) & (mul_34_17_n_11609 | mul_34_17_n_1961));
 assign mul_34_17_n_3553 = ((mul_34_17_n_1755 & mul_34_17_n_2447) | (mul_34_17_n_2898 & mul_34_17_n_2000));
 assign mul_34_17_n_3551 = ((mul_34_17_n_672 | mul_34_17_n_1059) & (mul_34_17_n_11552 | mul_34_17_n_1041));
 assign mul_34_17_n_3550 = ((mul_34_17_n_1754 | mul_34_17_n_2040) & (mul_34_17_n_11585 | mul_34_17_n_2681));
 assign mul_34_17_n_3549 = ((mul_34_17_n_674 | mul_34_17_n_1006) & (mul_34_17_n_11549 | mul_34_17_n_1005));
 assign mul_34_17_n_3548 = ~((mul_34_17_n_655 & mul_34_17_n_1648) | (mul_34_17_n_2902 & mul_34_17_n_1650));
 assign mul_34_17_n_3547 = ((mul_34_17_n_668 | mul_34_17_n_1174) & (mul_34_17_n_11558 | mul_34_17_n_1173));
 assign mul_34_17_n_3546 = ~((mul_34_17_n_1757 & mul_34_17_n_1774) | (mul_34_17_n_2900 & mul_34_17_n_1668));
 assign mul_34_17_n_3544 = ~((mul_34_17_n_659 & mul_34_17_n_1482) | (mul_34_17_n_2906 & mul_34_17_n_1456));
 assign mul_34_17_n_3542 = ~((mul_34_17_n_1743 & mul_34_17_n_2505) | (mul_34_17_n_2882 & mul_34_17_n_1880));
 assign mul_34_17_n_3541 = ((mul_34_17_n_1756 | mul_34_17_n_1768) & (mul_34_17_n_11582 | mul_34_17_n_1673));
 assign mul_34_17_n_3539 = ~((mul_34_17_n_657 & mul_34_17_n_1550) | (mul_34_17_n_2904 & mul_34_17_n_1555));
 assign mul_34_17_n_3538 = ((mul_34_17_n_1754 | mul_34_17_n_2083) & (mul_34_17_n_11585 | mul_34_17_n_1906));
 assign mul_34_17_n_3537 = ((mul_34_17_n_664 | mul_34_17_n_1300) & (mul_34_17_n_11564 | mul_34_17_n_1262));
 assign mul_34_17_n_3536 = ((mul_34_17_n_1744 | mul_34_17_n_2204) & (mul_34_17_n_11600 | mul_34_17_n_1917));
 assign mul_34_17_n_3534 = ~((mul_34_17_n_1735 & mul_34_17_n_2591) | (mul_34_17_n_2896 & mul_34_17_n_2323));
 assign mul_34_17_n_3533 = ((mul_34_17_n_1754 | mul_34_17_n_1921) & (mul_34_17_n_11585 | mul_34_17_n_2005));
 assign mul_34_17_n_3531 = ((mul_34_17_n_1734 | mul_34_17_n_2186) & (mul_34_17_n_11588 | mul_34_17_n_2315));
 assign mul_34_17_n_3530 = ((mul_34_17_n_1736 | mul_34_17_n_2652) & (mul_34_17_n_11591 | mul_34_17_n_2001));
 assign mul_34_17_n_3529 = ~((mul_34_17_n_665 & mul_34_17_n_1258) | (mul_34_17_n_2912 & mul_34_17_n_1301));
 assign mul_34_17_n_3527 = ((mul_34_17_n_1736 | mul_34_17_n_2207) & (mul_34_17_n_11591 | mul_34_17_n_2206));
 assign mul_34_17_n_3526 = ~((mul_34_17_n_687 & mul_34_17_n_711) | (mul_34_17_n_2933 & mul_34_17_n_712));
 assign mul_34_17_n_3525 = ((mul_34_17_n_1754 | mul_34_17_n_2078) & (mul_34_17_n_11585 | mul_34_17_n_2478));
 assign mul_34_17_n_3523 = ~((mul_34_17_n_1747 & mul_34_17_n_2570) | (mul_34_17_n_11593 & mul_34_17_n_2116));
 assign mul_34_17_n_3522 = ~((mul_34_17_n_655 & mul_34_17_n_1620) | (mul_34_17_n_2902 & mul_34_17_n_1639));
 assign mul_34_17_n_3521 = ~((mul_34_17_n_659 & mul_34_17_n_1470) | (mul_34_17_n_2906 & mul_34_17_n_1472));
 assign mul_34_17_n_3520 = ~((mul_34_17_n_1745 & mul_34_17_n_2561) | (mul_34_17_n_2888 & mul_34_17_n_2340));
 assign mul_34_17_n_3519 = ((mul_34_17_n_682 | mul_34_17_n_636) & (mul_34_17_n_11537 | mul_34_17_n_831));
 assign mul_34_17_n_3518 = ~((mul_34_17_n_1757 & mul_34_17_n_1773) | (mul_34_17_n_2900 & mul_34_17_n_955));
 assign mul_34_17_n_3517 = ~((mul_34_17_n_1745 & mul_34_17_n_2072) | (mul_34_17_n_2888 & mul_34_17_n_2175));
 assign mul_34_17_n_3516 = ~((mul_34_17_n_1751 & mul_34_17_n_2064) | (mul_34_17_n_2880 & mul_34_17_n_2063));
 assign mul_34_17_n_3515 = ~((mul_34_17_n_1739 & mul_34_17_n_2209) | (mul_34_17_n_2884 & mul_34_17_n_2123));
 assign mul_34_17_n_3513 = ~((mul_34_17_n_1745 & mul_34_17_n_2138) | (mul_34_17_n_2888 & mul_34_17_n_2016));
 assign mul_34_17_n_3512 = ((mul_34_17_n_657 & mul_34_17_n_1571) | (mul_34_17_n_2904 & mul_34_17_n_1572));
 assign mul_34_17_n_3511 = ((mul_34_17_n_654 | mul_34_17_n_1598) & (mul_34_17_n_11579 | mul_34_17_n_1627));
 assign mul_34_17_n_3510 = ((mul_34_17_n_1734 | mul_34_17_n_2368) & (mul_34_17_n_11588 | mul_34_17_n_2701));
 assign mul_34_17_n_3509 = ((mul_34_17_n_1740 | mul_34_17_n_2216) & (mul_34_17_n_11603 | mul_34_17_n_2322));
 assign mul_34_17_n_3508 = ((mul_34_17_n_657 & mul_34_17_n_1573) | (mul_34_17_n_2904 & mul_34_17_n_1540));
 assign mul_34_17_n_3507 = ((mul_34_17_n_1754 | mul_34_17_n_2495) & (mul_34_17_n_11585 | mul_34_17_n_1981));
 assign mul_34_17_n_3506 = ~((mul_34_17_n_1747 & mul_34_17_n_2007) | (mul_34_17_n_11593 & mul_34_17_n_2299));
 assign mul_34_17_n_3505 = ((mul_34_17_n_1757 & mul_34_17_n_1414) | (mul_34_17_n_2900 & mul_34_17_n_1111));
 assign mul_34_17_n_3503 = ((mul_34_17_n_1756 | mul_34_17_n_1758) & (mul_34_17_n_11582 | mul_34_17_n_1672));
 assign mul_34_17_n_3501 = ((mul_34_17_n_1736 | mul_34_17_n_2419) & (mul_34_17_n_11591 | mul_34_17_n_2525));
 assign mul_34_17_n_3500 = ((mul_34_17_n_655 & mul_34_17_n_1618) | (mul_34_17_n_2902 & mul_34_17_n_1633));
 assign mul_34_17_n_3499 = ~((mul_34_17_n_661 & mul_34_17_n_1429) | (mul_34_17_n_2908 & mul_34_17_n_1388));
 assign mul_34_17_n_3497 = ~((mul_34_17_n_681 & mul_34_17_n_838) | (mul_34_17_n_2928 & mul_34_17_n_853));
 assign mul_34_17_n_3496 = ((mul_34_17_n_1750 | mul_34_17_n_2448) & (mul_34_17_n_11612 | mul_34_17_n_2508));
 assign mul_34_17_n_3494 = ((mul_34_17_n_658 | mul_34_17_n_1449) & (mul_34_17_n_11573 | mul_34_17_n_1469));
 assign mul_34_17_n_3493 = ((mul_34_17_n_660 | mul_34_17_n_1395) & (mul_34_17_n_11570 | mul_34_17_n_1376));
 assign mul_34_17_n_3492 = ((mul_34_17_n_1737 & mul_34_17_n_2223) | (mul_34_17_n_2894 & mul_34_17_n_2221));
 assign mul_34_17_n_3491 = ~((mul_34_17_n_671 & mul_34_17_n_1117) | (mul_34_17_n_2918 & mul_34_17_n_1110));
 assign mul_34_17_n_3490 = ((mul_34_17_n_668 | mul_34_17_n_1127) & (mul_34_17_n_11558 | mul_34_17_n_1181));
 assign mul_34_17_n_3489 = ((mul_34_17_n_1754 | mul_34_17_n_1999) & (mul_34_17_n_11585 | mul_34_17_n_2628));
 assign mul_34_17_n_3488 = ~((mul_34_17_n_1747 & mul_34_17_n_2366) | (mul_34_17_n_11593 & mul_34_17_n_2638));
 assign mul_34_17_n_3487 = ((mul_34_17_n_664 | mul_34_17_n_1303) & (mul_34_17_n_11564 | mul_34_17_n_1300));
 assign mul_34_17_n_3486 = ~((mul_34_17_n_657 & mul_34_17_n_1558) | (mul_34_17_n_2904 & mul_34_17_n_1584));
 assign mul_34_17_n_3485 = ((mul_34_17_n_1746 | mul_34_17_n_2519) & (mul_34_17_n_11660 | mul_34_17_n_2003));
 assign mul_34_17_n_3484 = ((mul_34_17_n_1738 | mul_34_17_n_1927) & (mul_34_17_n_11606 | mul_34_17_n_2372));
 assign mul_34_17_n_3483 = ~((mul_34_17_n_663 & mul_34_17_n_1340) | (mul_34_17_n_2910 & mul_34_17_n_1318));
 assign mul_34_17_n_3482 = ((mul_34_17_n_1746 | mul_34_17_n_2280) & (mul_34_17_n_11672 | mul_34_17_n_2696));
 assign mul_34_17_n_3481 = ((mul_34_17_n_686 | mul_34_17_n_714) & (mul_34_17_n_11531 | mul_34_17_n_722));
 assign mul_34_17_n_3480 = ~((mul_34_17_n_685 & mul_34_17_n_773) | (mul_34_17_n_2931 & mul_34_17_n_800));
 assign mul_34_17_n_3479 = ((mul_34_17_n_656 | mul_34_17_n_1539) & (mul_34_17_n_11576 | mul_34_17_n_1544));
 assign mul_34_17_n_3478 = ~((mul_34_17_n_1741 & mul_34_17_n_2451) | (mul_34_17_n_2886 & mul_34_17_n_1868));
 assign mul_34_17_n_3477 = ~((mul_34_17_n_1755 & mul_34_17_n_2668) | (mul_34_17_n_2898 & mul_34_17_n_2170));
 assign mul_34_17_n_3476 = ((mul_34_17_n_1752 | mul_34_17_n_2091) & (mul_34_17_n_11615 | mul_34_17_n_2410));
 assign mul_34_17_n_3475 = ((mul_34_17_n_1740 | mul_34_17_n_1902) & (mul_34_17_n_11603 | mul_34_17_n_2038));
 assign mul_34_17_n_3474 = ~((mul_34_17_n_1751 & mul_34_17_n_2459) | (mul_34_17_n_2880 & mul_34_17_n_2050));
 assign mul_34_17_n_3473 = ~((mul_34_17_n_687 & mul_34_17_n_807) | (mul_34_17_n_2933 & mul_34_17_n_707));
 assign mul_34_17_n_3472 = ~((mul_34_17_n_1739 & mul_34_17_n_2195) | (mul_34_17_n_2884 & mul_34_17_n_2579));
 assign mul_34_17_n_3471 = ~((mul_34_17_n_1751 & mul_34_17_n_1987) | (mul_34_17_n_2880 & mul_34_17_n_2047));
 assign mul_34_17_n_3470 = ((mul_34_17_n_656 | mul_34_17_n_1581) & (mul_34_17_n_11576 | mul_34_17_n_1522));
 assign mul_34_17_n_3469 = ~((mul_34_17_n_1735 & mul_34_17_n_2455) | (mul_34_17_n_2896 & mul_34_17_n_2127));
 assign mul_34_17_n_3468 = ~((mul_34_17_n_1739 & mul_34_17_n_2586) | (mul_34_17_n_2884 & mul_34_17_n_2046));
 assign mul_34_17_n_3467 = ~((mul_34_17_n_1749 & mul_34_17_n_2101) | (mul_34_17_n_2890 & mul_34_17_n_2337));
 assign mul_34_17_n_3466 = ((mul_34_17_n_1742 | mul_34_17_n_1851) & (mul_34_17_n_11609 | mul_34_17_n_2102));
 assign mul_34_17_n_3465 = ~((mul_34_17_n_691 & mul_34_17_n_1009) | (mul_34_17_n_2936 & mul_34_17_n_705));
 assign mul_34_17_n_3464 = ~((mul_34_17_n_661 & mul_34_17_n_1435) | (mul_34_17_n_2908 & mul_34_17_n_1386));
 assign mul_34_17_n_3463 = ~((mul_34_17_n_1749 & mul_34_17_n_1890) | (mul_34_17_n_2890 & mul_34_17_n_2044));
 assign mul_34_17_n_3462 = ((mul_34_17_n_688 | mul_34_17_n_731) & (mul_34_17_n_11528 | mul_34_17_n_696));
 assign mul_34_17_n_3461 = ((mul_34_17_n_1744 | mul_34_17_n_2693) & (mul_34_17_n_11600 | mul_34_17_n_2176));
 assign mul_34_17_n_3460 = ~((mul_34_17_n_661 & mul_34_17_n_1439) | (mul_34_17_n_2908 & mul_34_17_n_1396));
 assign mul_34_17_n_3459 = ~((mul_34_17_n_1743 & mul_34_17_n_2454) | (mul_34_17_n_2882 & mul_34_17_n_2384));
 assign mul_34_17_n_3458 = ~((mul_34_17_n_1749 & mul_34_17_n_1905) | (mul_34_17_n_2890 & mul_34_17_n_2039));
 assign mul_34_17_n_3457 = ((mul_34_17_n_674 | mul_34_17_n_978) & (mul_34_17_n_11549 | mul_34_17_n_1004));
 assign mul_34_17_n_3456 = ((mul_34_17_n_658 | mul_34_17_n_1485) & (mul_34_17_n_11573 | mul_34_17_n_1488));
 assign mul_34_17_n_3455 = ((mul_34_17_n_1744 | mul_34_17_n_2474) & (mul_34_17_n_11600 | mul_34_17_n_2480));
 assign mul_34_17_n_3454 = ((mul_34_17_n_1738 | mul_34_17_n_2504) & (mul_34_17_n_11606 | mul_34_17_n_2499));
 assign mul_34_17_n_3453 = ((mul_34_17_n_654 | mul_34_17_n_1631) & (mul_34_17_n_11579 | mul_34_17_n_1596));
 assign mul_34_17_n_3452 = ((mul_34_17_n_1736 | mul_34_17_n_2407) & (mul_34_17_n_11591 | mul_34_17_n_2037));
 assign mul_34_17_n_3451 = ~((mul_34_17_n_1737 & mul_34_17_n_2427) | (mul_34_17_n_2894 & mul_34_17_n_2355));
 assign mul_34_17_n_3450 = ((mul_34_17_n_670 | mul_34_17_n_1123) & (mul_34_17_n_11555 | mul_34_17_n_1090));
 assign mul_34_17_n_3449 = ((mul_34_17_n_662 | mul_34_17_n_1358) & (mul_34_17_n_11567 | mul_34_17_n_1348));
 assign mul_34_17_n_3448 = ((mul_34_17_n_1742 | mul_34_17_n_2183) & (mul_34_17_n_11609 | mul_34_17_n_2348));
 assign mul_34_17_n_3447 = ((mul_34_17_n_666 | mul_34_17_n_1213) & (mul_34_17_n_11561 | mul_34_17_n_1234));
 assign mul_34_17_n_3446 = ((mul_34_17_n_668 | mul_34_17_n_1128) & (mul_34_17_n_11558 | mul_34_17_n_1172));
 assign mul_34_17_n_3445 = ~((mul_34_17_n_1749 & mul_34_17_n_2369) | (mul_34_17_n_2890 & mul_34_17_n_1899));
 assign mul_34_17_n_3444 = ((mul_34_17_n_688 | mul_34_17_n_697) & (mul_34_17_n_11528 | mul_34_17_n_708));
 assign mul_34_17_n_3442 = ((mul_34_17_n_1746 | mul_34_17_n_2320) & (mul_34_17_n_11646 | mul_34_17_n_2184));
 assign mul_34_17_n_3441 = ~((mul_34_17_n_1755 & mul_34_17_n_1982) | (mul_34_17_n_2898 & mul_34_17_n_2452));
 assign mul_34_17_n_3440 = ~((mul_34_17_n_1753 & mul_34_17_n_1978) | (mul_34_17_n_2878 & mul_34_17_n_2192));
 assign mul_34_17_n_3439 = ((mul_34_17_n_654 | mul_34_17_n_1611) & (mul_34_17_n_11579 | mul_34_17_n_1600));
 assign mul_34_17_n_3438 = ((mul_34_17_n_684 | mul_34_17_n_770) & (mul_34_17_n_11534 | mul_34_17_n_763));
 assign mul_34_17_n_3437 = ~((mul_34_17_n_1740 | mul_34_17_n_1859) & (mul_34_17_n_11603 | mul_34_17_n_2158));
 assign mul_34_17_n_3436 = ~((mul_34_17_n_656 | mul_34_17_n_1544) & (mul_34_17_n_11576 | mul_34_17_n_1562));
 assign mul_34_17_n_3435 = ((mul_34_17_n_1736 | mul_34_17_n_1887) & (mul_34_17_n_11591 | mul_34_17_n_2419));
 assign mul_34_17_n_3434 = ~((mul_34_17_n_654 | mul_34_17_n_1596) & (mul_34_17_n_11579 | mul_34_17_n_1651));
 assign mul_34_17_n_3433 = ((mul_34_17_n_672 | mul_34_17_n_1041) & (mul_34_17_n_11552 | mul_34_17_n_1023));
 assign mul_34_17_n_3432 = ~((mul_34_17_n_661 & mul_34_17_n_1386) | (mul_34_17_n_2908 & mul_34_17_n_1438));
 assign mul_34_17_n_3431 = ((mul_34_17_n_1734 | mul_34_17_n_2494) & (mul_34_17_n_11588 | mul_34_17_n_2234));
 assign mul_34_17_n_3430 = ((mul_34_17_n_1736 | mul_34_17_n_2037) & (mul_34_17_n_11591 | mul_34_17_n_2674));
 assign mul_34_17_n_3429 = ((mul_34_17_n_682 | mul_34_17_n_804) & (mul_34_17_n_11537 | mul_34_17_n_810));
 assign mul_34_17_n_3428 = ~((mul_34_17_n_671 & mul_34_17_n_1072) | (mul_34_17_n_2918 & mul_34_17_n_1101));
 assign mul_34_17_n_3427 = ((mul_34_17_n_676 | mul_34_17_n_926) & (mul_34_17_n_11546 | mul_34_17_n_921));
 assign mul_34_17_n_3426 = ~((mul_34_17_n_685 & mul_34_17_n_787) | (mul_34_17_n_2931 & mul_34_17_n_790));
 assign mul_34_17_n_3425 = ((mul_34_17_n_1753 & mul_34_17_n_2622) | (mul_34_17_n_2878 & mul_34_17_n_2021));
 assign mul_34_17_n_3424 = ((mul_34_17_n_664 | mul_34_17_n_1273) & (mul_34_17_n_11564 | mul_34_17_n_1303));
 assign mul_34_17_n_3423 = ~((mul_34_17_n_1734 | mul_34_17_n_2173) & (mul_34_17_n_11588 | mul_34_17_n_2171));
 assign mul_34_17_n_3422 = ((mul_34_17_n_1738 | mul_34_17_n_2571) & (mul_34_17_n_11606 | mul_34_17_n_2053));
 assign mul_34_17_n_3421 = ((mul_34_17_n_1740 | mul_34_17_n_2231) & (mul_34_17_n_11603 | mul_34_17_n_2236));
 assign mul_34_17_n_3420 = ((mul_34_17_n_686 | mul_34_17_n_730) & (mul_34_17_n_11531 | mul_34_17_n_713));
 assign mul_34_17_n_3419 = ((mul_34_17_n_676 | mul_34_17_n_947) & (mul_34_17_n_11546 | mul_34_17_n_920));
 assign mul_34_17_n_3418 = ((mul_34_17_n_671 & mul_34_17_n_1070) | (mul_34_17_n_2918 & mul_34_17_n_1106));
 assign mul_34_17_n_3417 = ((mul_34_17_n_1756 | mul_34_17_n_903) & (mul_34_17_n_11582 | mul_34_17_n_1772));
 assign mul_34_17_n_3415 = ((mul_34_17_n_1740 | mul_34_17_n_1867) & (mul_34_17_n_11603 | mul_34_17_n_2093));
 assign mul_34_17_n_3414 = ((mul_34_17_n_668 | mul_34_17_n_1159) & (mul_34_17_n_11558 | mul_34_17_n_1131));
 assign mul_34_17_n_3413 = ~((mul_34_17_n_1754 | mul_34_17_n_2628) & (mul_34_17_n_11585 | mul_34_17_n_2610));
 assign mul_34_17_n_3412 = ~((mul_34_17_n_1750 | mul_34_17_n_2051) & (mul_34_17_n_11612 | mul_34_17_n_2129));
 assign mul_34_17_n_3411 = ((mul_34_17_n_1756 | mul_34_17_n_1670) & (mul_34_17_n_11582 | mul_34_17_n_1687));
 assign mul_34_17_n_3410 = ((mul_34_17_n_666 | mul_34_17_n_1226) & (mul_34_17_n_11561 | mul_34_17_n_1215));
 assign mul_34_17_n_3409 = ~((mul_34_17_n_674 | mul_34_17_n_970) & (mul_34_17_n_11549 | mul_34_17_n_980));
 assign mul_34_17_n_3408 = ~((mul_34_17_n_1734 | mul_34_17_n_2128) & (mul_34_17_n_11588 | mul_34_17_n_2607));
 assign mul_34_17_n_3407 = ((mul_34_17_n_1738 | mul_34_17_n_2499) & (mul_34_17_n_11606 | mul_34_17_n_2351));
 assign mul_34_17_n_3406 = ((mul_34_17_n_1750 | mul_34_17_n_1692) & (mul_34_17_n_11612 | mul_34_17_n_2067));
 assign mul_34_17_n_3405 = ~((mul_34_17_n_685 & mul_34_17_n_781) | (mul_34_17_n_2931 & mul_34_17_n_798));
 assign mul_34_17_n_3403 = ((mul_34_17_n_1734 | mul_34_17_n_2646) & (mul_34_17_n_11588 | mul_34_17_n_2414));
 assign mul_34_17_n_3402 = ((mul_34_17_n_1756 | mul_34_17_n_2614) & (mul_34_17_n_11582 | mul_34_17_n_2256));
 assign mul_34_17_n_3401 = ~((mul_34_17_n_1757 & mul_34_17_n_1975) | (mul_34_17_n_2900 & mul_34_17_n_2435));
 assign mul_34_17_n_3399 = ((mul_34_17_n_664 | mul_34_17_n_1254) & (mul_34_17_n_11564 | mul_34_17_n_1304));
 assign mul_34_17_n_3397 = ((mul_34_17_n_1738 | mul_34_17_n_2110) & (mul_34_17_n_11606 | mul_34_17_n_1854));
 assign mul_34_17_n_3395 = ((mul_34_17_n_1740 | mul_34_17_n_2336) & (mul_34_17_n_11603 | mul_34_17_n_1902));
 assign mul_34_17_n_3393 = ((mul_34_17_n_1750 | mul_34_17_n_2640) & (mul_34_17_n_11612 | mul_34_17_n_1986));
 assign mul_34_17_n_3391 = ~((mul_34_17_n_654 | mul_34_17_n_1612) & (mul_34_17_n_11579 | mul_34_17_n_1599));
 assign mul_34_17_n_3389 = ((mul_34_17_n_662 | mul_34_17_n_1317) & (mul_34_17_n_11567 | mul_34_17_n_1355));
 assign mul_34_17_n_3387 = ((mul_34_17_n_1742 | mul_34_17_n_2383) & (mul_34_17_n_11609 | mul_34_17_n_2634));
 assign mul_34_17_n_3386 = ((mul_34_17_n_660 | mul_34_17_n_1407) & (mul_34_17_n_11570 | mul_34_17_n_1392));
 assign mul_34_17_n_3385 = ((mul_34_17_n_1752 | mul_34_17_n_2262) & (mul_34_17_n_11615 | mul_34_17_n_2107));
 assign mul_34_17_n_3384 = ~((mul_34_17_n_1756 | mul_34_17_n_1775) & (mul_34_17_n_11582 | mul_34_17_n_1669));
 assign mul_34_17_n_3383 = ~((mul_34_17_n_1738 | mul_34_17_n_2045) & (mul_34_17_n_11606 | mul_34_17_n_2098));
 assign mul_34_17_n_3382 = ((mul_34_17_n_654 | mul_34_17_n_1652) & (mul_34_17_n_11579 | mul_34_17_n_1603));
 assign mul_34_17_n_3381 = ((mul_34_17_n_1742 | mul_34_17_n_2102) & (mul_34_17_n_11609 | mul_34_17_n_2592));
 assign mul_34_17_n_3380 = ((mul_34_17_n_1734 | mul_34_17_n_2167) & (mul_34_17_n_11588 | mul_34_17_n_2075));
 assign mul_34_17_n_3379 = ((mul_34_17_n_656 | mul_34_17_n_1536) & (mul_34_17_n_11576 | mul_34_17_n_1579));
 assign mul_34_17_n_3378 = ~((mul_34_17_n_664 | mul_34_17_n_1260) & (mul_34_17_n_11564 | mul_34_17_n_1267));
 assign mul_34_17_n_3377 = ((mul_34_17_n_654 | mul_34_17_n_1600) & (mul_34_17_n_11579 | mul_34_17_n_1598));
 assign mul_34_17_n_3376 = ((mul_34_17_n_1734 | mul_34_17_n_2234) & (mul_34_17_n_11588 | mul_34_17_n_2049));
 assign mul_34_17_n_3375 = ((mul_34_17_n_678 | mul_34_17_n_876) & (mul_34_17_n_11543 | mul_34_17_n_917));
 assign mul_34_17_n_3374 = ~((mul_34_17_n_1741 & mul_34_17_n_2589) | (mul_34_17_n_2886 & mul_34_17_n_1853));
 assign mul_34_17_n_3373 = ~((mul_34_17_n_1747 & mul_34_17_n_2212) | (mul_34_17_n_11593 & mul_34_17_n_2226));
 assign mul_34_17_n_3372 = ((mul_34_17_n_660 | mul_34_17_n_1398) & (mul_34_17_n_11570 | mul_34_17_n_1440));
 assign mul_34_17_n_3371 = ((mul_34_17_n_656 | mul_34_17_n_1570) & (mul_34_17_n_11576 | mul_34_17_n_1531));
 assign mul_34_17_n_3370 = ~((mul_34_17_n_1757 & mul_34_17_n_1175) | (mul_34_17_n_2900 & mul_34_17_n_2542));
 assign mul_34_17_n_3368 = ((mul_34_17_n_1742 | mul_34_17_n_2214) & (mul_34_17_n_11609 | mul_34_17_n_2160));
 assign mul_34_17_n_3367 = ((mul_34_17_n_656 | mul_34_17_n_1566) & (mul_34_17_n_11576 | mul_34_17_n_1557));
 assign mul_34_17_n_3366 = ~((mul_34_17_n_1757 & mul_34_17_n_1831) | (mul_34_17_n_2900 & mul_34_17_n_1414));
 assign mul_34_17_n_3365 = ~((mul_34_17_n_667 & mul_34_17_n_1206) | (mul_34_17_n_2914 & mul_34_17_n_1237));
 assign mul_34_17_n_3364 = ~((mul_34_17_n_657 & mul_34_17_n_1523) | (mul_34_17_n_2904 & mul_34_17_n_1520));
 assign mul_34_17_n_3363 = ((mul_34_17_n_688 | mul_34_17_n_708) & (mul_34_17_n_11528 | mul_34_17_n_731));
 assign mul_34_17_n_3362 = ((mul_34_17_n_1746 | mul_34_17_n_2663) & (mul_34_17_n_11682 | mul_34_17_n_2466));
 assign mul_34_17_n_3361 = ~((mul_34_17_n_677 & mul_34_17_n_944) | (mul_34_17_n_2924 & mul_34_17_n_935));
 assign mul_34_17_n_3360 = ~((mul_34_17_n_671 & mul_34_17_n_1098) | (mul_34_17_n_2918 & mul_34_17_n_1087));
 assign mul_34_17_n_3359 = ((mul_34_17_n_660 | mul_34_17_n_1381) & (mul_34_17_n_11570 | mul_34_17_n_1378));
 assign mul_34_17_n_3358 = ((mul_34_17_n_672 | mul_34_17_n_1026) & (mul_34_17_n_11552 | mul_34_17_n_1059));
 assign mul_34_17_n_3357 = ~((mul_34_17_n_1745 & mul_34_17_n_1875) | (mul_34_17_n_2888 & mul_34_17_n_1968));
 assign mul_34_17_n_3356 = ((mul_34_17_n_1736 | mul_34_17_n_2206) & (mul_34_17_n_11591 | mul_34_17_n_2208));
 assign mul_34_17_n_3355 = ((mul_34_17_n_654 | mul_34_17_n_1616) & (mul_34_17_n_11579 | mul_34_17_n_1614));
 assign mul_34_17_n_3354 = ((mul_34_17_n_1742 | mul_34_17_n_2248) & (mul_34_17_n_11609 | mul_34_17_n_1851));
 assign mul_34_17_n_3353 = ~((mul_34_17_n_657 & mul_34_17_n_1538) | (mul_34_17_n_2904 & mul_34_17_n_1561));
 assign mul_34_17_n_3351 = ((mul_34_17_n_1748 | mul_34_17_n_2230) & (mul_34_17_n_11597 | mul_34_17_n_1883));
 assign mul_34_17_n_3349 = ~((mul_34_17_n_1743 & mul_34_17_n_2333) | (mul_34_17_n_2882 & mul_34_17_n_2321));
 assign mul_34_17_n_3348 = ((mul_34_17_n_1744 | mul_34_17_n_1917) & (mul_34_17_n_11600 | mul_34_17_n_2641));
 assign mul_34_17_n_3347 = ((mul_34_17_n_1752 | mul_34_17_n_1998) & (mul_34_17_n_11615 | mul_34_17_n_2042));
 assign mul_34_17_n_3346 = ((mul_34_17_n_664 | mul_34_17_n_1278) & (mul_34_17_n_11564 | mul_34_17_n_1288));
 assign mul_34_17_n_3345 = ((mul_34_17_n_1746 | mul_34_17_n_2003) & (mul_34_17_n_11666 | mul_34_17_n_1946));
 assign mul_34_17_n_3344 = ((mul_34_17_n_656 | mul_34_17_n_1530) & (mul_34_17_n_11576 | mul_34_17_n_1537));
 assign mul_34_17_n_3343 = ((mul_34_17_n_654 | mul_34_17_n_1649) & (mul_34_17_n_11579 | mul_34_17_n_1644));
 assign mul_34_17_n_3341 = ((mul_34_17_n_1746 | mul_34_17_n_2696) & (mul_34_17_n_11679 | mul_34_17_n_2335));
 assign mul_34_17_n_3340 = ((mul_34_17_n_686 | mul_34_17_n_704) & (mul_34_17_n_11531 | mul_34_17_n_714));
 assign mul_34_17_n_3339 = ((mul_34_17_n_678 | mul_34_17_n_878) & (mul_34_17_n_11543 | mul_34_17_n_895));
 assign mul_34_17_n_3338 = ((mul_34_17_n_678 | mul_34_17_n_893) & (mul_34_17_n_11543 | mul_34_17_n_886));
 assign mul_34_17_n_3336 = ((mul_34_17_n_1750 | mul_34_17_n_2603) & (mul_34_17_n_11612 | mul_34_17_n_2640));
 assign mul_34_17_n_3335 = ~((mul_34_17_n_1753 & mul_34_17_n_2470) | (mul_34_17_n_2878 & mul_34_17_n_2114));
 assign mul_34_17_n_3334 = ((mul_34_17_n_654 | mul_34_17_n_1615) & (mul_34_17_n_11579 | mul_34_17_n_1611));
 assign mul_34_17_n_3333 = ((mul_34_17_n_680 | mul_34_17_n_840) & (mul_34_17_n_11540 | mul_34_17_n_864));
 assign mul_34_17_n_3332 = ~((mul_34_17_n_1741 & mul_34_17_n_2484) | (mul_34_17_n_2886 & mul_34_17_n_2568));
 assign mul_34_17_n_3330 = ~((mul_34_17_n_1757 & mul_34_17_n_1760) | (mul_34_17_n_2900 & mul_34_17_n_1682));
 assign mul_34_17_n_3329 = ((mul_34_17_n_664 | mul_34_17_n_1275) & (mul_34_17_n_11564 | mul_34_17_n_1255));
 assign mul_34_17_n_3328 = ((mul_34_17_n_1734 | mul_34_17_n_2414) & (mul_34_17_n_11588 | mul_34_17_n_2692));
 assign mul_34_17_n_3327 = ((mul_34_17_n_668 | mul_34_17_n_1172) & (mul_34_17_n_11558 | mul_34_17_n_1170));
 assign mul_34_17_n_3326 = ~((mul_34_17_n_661 & mul_34_17_n_1422) | (mul_34_17_n_2908 & mul_34_17_n_1402));
 assign mul_34_17_n_3324 = ~((mul_34_17_n_1749 & mul_34_17_n_1992) | (mul_34_17_n_2890 & mul_34_17_n_2341));
 assign mul_34_17_n_3323 = ((mul_34_17_n_678 | mul_34_17_n_882) & (mul_34_17_n_11543 | mul_34_17_n_890));
 assign mul_34_17_n_3322 = ~((mul_34_17_n_1741 & mul_34_17_n_2141) | (mul_34_17_n_2886 & mul_34_17_n_2151));
 assign mul_34_17_n_3321 = ~((mul_34_17_n_655 & mul_34_17_n_1663) | (mul_34_17_n_2902 & mul_34_17_n_1623));
 assign mul_34_17_n_3320 = ~((mul_34_17_n_1745 & mul_34_17_n_2095) | (mul_34_17_n_2888 & mul_34_17_n_2274));
 assign mul_34_17_n_3319 = ~((mul_34_17_n_1753 & mul_34_17_n_2192) | (mul_34_17_n_2878 & mul_34_17_n_2590));
 assign mul_34_17_n_3317 = ~((mul_34_17_n_1751 & mul_34_17_n_2312) | (mul_34_17_n_2880 & mul_34_17_n_2043));
 assign mul_34_17_n_3316 = ((mul_34_17_n_1740 | mul_34_17_n_1952) & (mul_34_17_n_11603 | mul_34_17_n_1938));
 assign mul_34_17_n_3315 = ((mul_34_17_n_1734 | mul_34_17_n_1922) & (mul_34_17_n_11588 | mul_34_17_n_2633));
 assign mul_34_17_n_3314 = ~((mul_34_17_n_1739 & mul_34_17_n_1948) | (mul_34_17_n_2884 & mul_34_17_n_2187));
 assign mul_34_17_n_3313 = ((mul_34_17_n_662 | mul_34_17_n_1363) & (mul_34_17_n_11567 | mul_34_17_n_1321));
 assign mul_34_17_n_3311 = ~((mul_34_17_n_1741 & mul_34_17_n_2279) | (mul_34_17_n_2886 & mul_34_17_n_1973));
 assign mul_34_17_n_3310 = ((mul_34_17_n_1748 | mul_34_17_n_2111) & (mul_34_17_n_11597 | mul_34_17_n_2509));
 assign mul_34_17_n_3309 = ((mul_34_17_n_658 | mul_34_17_n_1496) & (mul_34_17_n_11573 | mul_34_17_n_1481));
 assign mul_34_17_n_3308 = ((mul_34_17_n_1752 | mul_34_17_n_2539) & (mul_34_17_n_11615 | mul_34_17_n_1983));
 assign mul_34_17_n_3307 = ~((mul_34_17_n_1747 & mul_34_17_n_1870) | (mul_34_17_n_11593 & mul_34_17_n_2153));
 assign mul_34_17_n_3306 = ((mul_34_17_n_668 | mul_34_17_n_1134) & (mul_34_17_n_11558 | mul_34_17_n_1156));
 assign mul_34_17_n_3305 = ~((mul_34_17_n_677 & mul_34_17_n_922) | (mul_34_17_n_2924 & mul_34_17_n_952));
 assign mul_34_17_n_3304 = ((mul_34_17_n_664 | mul_34_17_n_1276) & (mul_34_17_n_11564 | mul_34_17_n_1256));
 assign mul_34_17_n_3303 = ((mul_34_17_n_666 | mul_34_17_n_1227) & (mul_34_17_n_11561 | mul_34_17_n_1208));
 assign mul_34_17_n_3302 = ((mul_34_17_n_680 | mul_34_17_n_849) & (mul_34_17_n_11540 | mul_34_17_n_845));
 assign mul_34_17_n_3301 = ((mul_34_17_n_676 | mul_34_17_n_934) & (mul_34_17_n_11546 | mul_34_17_n_958));
 assign mul_34_17_n_3300 = ~((mul_34_17_n_657 & mul_34_17_n_1572) | (mul_34_17_n_2904 & mul_34_17_n_1548));
 assign mul_34_17_n_3299 = ((mul_34_17_n_1748 | mul_34_17_n_2374) & (mul_34_17_n_11597 | mul_34_17_n_2084));
 assign mul_34_17_n_3298 = ~((mul_34_17_n_663 & mul_34_17_n_1364) | (mul_34_17_n_2910 & mul_34_17_n_1344));
 assign mul_34_17_n_3297 = ((mul_34_17_n_1748 | mul_34_17_n_2645) & (mul_34_17_n_11597 | mul_34_17_n_2574));
 assign mul_34_17_n_3296 = ~((mul_34_17_n_654 | mul_34_17_n_1659) & (mul_34_17_n_11579 | mul_34_17_n_1617));
 assign mul_34_17_n_3295 = ((mul_34_17_n_1736 | mul_34_17_n_2181) & (mul_34_17_n_11591 | mul_34_17_n_2436));
 assign mul_34_17_n_3294 = ~((mul_34_17_n_1751 & mul_34_17_n_2679) | (mul_34_17_n_2880 & mul_34_17_n_2635));
 assign mul_34_17_n_3293 = ~((mul_34_17_n_1739 & mul_34_17_n_2203) | (mul_34_17_n_2884 & mul_34_17_n_1934));
 assign mul_34_17_n_3291 = ((mul_34_17_n_1734 | mul_34_17_n_1912) & (mul_34_17_n_11588 | mul_34_17_n_2194));
 assign mul_34_17_n_3289 = ((mul_34_17_n_1754 | mul_34_17_n_1937) & (mul_34_17_n_11585 | mul_34_17_n_2608));
 assign mul_34_17_n_3288 = ((mul_34_17_n_1746 | mul_34_17_n_2117) & (mul_34_17_n_11658 | mul_34_17_n_1935));
 assign mul_34_17_n_3287 = ((mul_34_17_n_658 | mul_34_17_n_1491) & (mul_34_17_n_11573 | mul_34_17_n_1471));
 assign mul_34_17_n_3286 = ~((mul_34_17_n_1747 & mul_34_17_n_2299) | (mul_34_17_n_11593 & mul_34_17_n_1931));
 assign mul_34_17_n_3285 = ~((mul_34_17_n_1745 & mul_34_17_n_2273) | (mul_34_17_n_2888 & mul_34_17_n_2228));
 assign mul_34_17_n_3284 = ~((mul_34_17_n_1736 | mul_34_17_n_1932) & (mul_34_17_n_11591 | mul_34_17_n_2215));
 assign mul_34_17_n_3283 = ~((mul_34_17_n_1756 | mul_34_17_n_1770) & (mul_34_17_n_11582 | mul_34_17_n_1670));
 assign mul_34_17_n_3282 = ((mul_34_17_n_660 | mul_34_17_n_1443) & (mul_34_17_n_11570 | mul_34_17_n_1389));
 assign mul_34_17_n_3281 = ((mul_34_17_n_672 | mul_34_17_n_1042) & (mul_34_17_n_11552 | mul_34_17_n_1045));
 assign mul_34_17_n_3280 = ((mul_34_17_n_1746 | mul_34_17_n_2297) & (mul_34_17_n_11651 | mul_34_17_n_2189));
 assign mul_34_17_n_3279 = ((mul_34_17_n_672 | mul_34_17_n_1017) & (mul_34_17_n_11552 | mul_34_17_n_1048));
 assign mul_34_17_n_3278 = ((mul_34_17_n_686 | mul_34_17_n_722) & (mul_34_17_n_11531 | mul_34_17_n_730));
 assign mul_34_17_n_3277 = ((mul_34_17_n_662 | mul_34_17_n_1370) & (mul_34_17_n_11567 | mul_34_17_n_1349));
 assign mul_34_17_n_3276 = ((mul_34_17_n_654 | mul_34_17_n_1594) & (mul_34_17_n_11579 | mul_34_17_n_1643));
 assign mul_34_17_n_3275 = ~((mul_34_17_n_669 & mul_34_17_n_1177) | (mul_34_17_n_2916 & mul_34_17_n_1126));
 assign mul_34_17_n_3274 = ((mul_34_17_n_662 | mul_34_17_n_1368) & (mul_34_17_n_11567 | mul_34_17_n_1363));
 assign mul_34_17_n_3273 = ((mul_34_17_n_658 | mul_34_17_n_1481) & (mul_34_17_n_11573 | mul_34_17_n_1461));
 assign mul_34_17_n_3271 = ~((mul_34_17_n_655 & mul_34_17_n_1593) | (mul_34_17_n_2902 & mul_34_17_n_1624));
 assign mul_34_17_n_3269 = ((mul_34_17_n_656 | mul_34_17_n_1529) & (mul_34_17_n_11576 | mul_34_17_n_1524));
 assign mul_34_17_n_3267 = ((mul_34_17_n_1748 | mul_34_17_n_2084) & (mul_34_17_n_11597 | mul_34_17_n_2302));
 assign mul_34_17_n_3266 = ((mul_34_17_n_662 | mul_34_17_n_1349) & (mul_34_17_n_11567 | mul_34_17_n_1327));
 assign mul_34_17_n_3265 = ((mul_34_17_n_1752 | mul_34_17_n_1929) & (mul_34_17_n_11615 | mul_34_17_n_1998));
 assign mul_34_17_n_3264 = ((mul_34_17_n_660 | mul_34_17_n_1417) & (mul_34_17_n_11570 | mul_34_17_n_1420));
 assign mul_34_17_n_3263 = ((mul_34_17_n_666 | mul_34_17_n_1235) & (mul_34_17_n_11561 | mul_34_17_n_1185));
 assign mul_34_17_n_3262 = ((mul_34_17_n_688 | mul_34_17_n_698) & (mul_34_17_n_11528 | mul_34_17_n_697));
 assign mul_34_17_n_3261 = ~((mul_34_17_n_655 & mul_34_17_n_1606) | (mul_34_17_n_2902 & mul_34_17_n_1628));
 assign mul_34_17_n_3259 = ~((mul_34_17_n_1749 & mul_34_17_n_2011) | (mul_34_17_n_2890 & mul_34_17_n_2210));
 assign mul_34_17_n_3258 = ((mul_34_17_n_672 | mul_34_17_n_1027) & (mul_34_17_n_11552 | mul_34_17_n_1024));
 assign mul_34_17_n_3257 = ~((mul_34_17_n_659 & mul_34_17_n_1507) | (mul_34_17_n_2906 & mul_34_17_n_1479));
 assign mul_34_17_n_3256 = ~((mul_34_17_n_1737 & mul_34_17_n_2503) | (mul_34_17_n_2894 & mul_34_17_n_2245));
 assign mul_34_17_n_3255 = ((mul_34_17_n_654 | mul_34_17_n_1644) & (mul_34_17_n_11579 | mul_34_17_n_1590));
 assign mul_34_17_n_3254 = ((mul_34_17_n_1738 | mul_34_17_n_2052) & (mul_34_17_n_11606 | mul_34_17_n_1927));
 assign mul_34_17_n_3253 = ((mul_34_17_n_676 | mul_34_17_n_949) & (mul_34_17_n_11546 | mul_34_17_n_956));
 assign mul_34_17_n_3252 = ((mul_34_17_n_666 | mul_34_17_n_1230) & (mul_34_17_n_11561 | mul_34_17_n_1196));
 assign mul_34_17_n_3251 = ((mul_34_17_n_1738 | mul_34_17_n_2125) & (mul_34_17_n_11606 | mul_34_17_n_2685));
 assign mul_34_17_n_3250 = ~((mul_34_17_n_1735 & mul_34_17_n_2521) | (mul_34_17_n_2896 & mul_34_17_n_2565));
 assign mul_34_17_n_3249 = ((mul_34_17_n_1754 | mul_34_17_n_1916) & (mul_34_17_n_11585 | mul_34_17_n_2083));
 assign mul_34_17_n_3248 = ((mul_34_17_n_658 | mul_34_17_n_1478) & (mul_34_17_n_11573 | mul_34_17_n_1473));
 assign mul_34_17_n_3246 = ((mul_34_17_n_1744 | mul_34_17_n_2329) & (mul_34_17_n_11600 | mul_34_17_n_2204));
 assign mul_34_17_n_3244 = ((mul_34_17_n_668 | mul_34_17_n_1149) & (mul_34_17_n_11558 | mul_34_17_n_1162));
 assign mul_34_17_n_3243 = ((mul_34_17_n_674 | mul_34_17_n_999) & (mul_34_17_n_11549 | mul_34_17_n_1006));
 assign mul_34_17_n_3241 = ((mul_34_17_n_1750 | mul_34_17_n_2531) & (mul_34_17_n_11612 | mul_34_17_n_2019));
 assign mul_34_17_n_3239 = ((mul_34_17_n_1748 | mul_34_17_n_2538) & (mul_34_17_n_11597 | mul_34_17_n_2029));
 assign mul_34_17_n_3238 = ~((mul_34_17_n_1736 | mul_34_17_n_2523) & (mul_34_17_n_11591 | mul_34_17_n_2407));
 assign mul_34_17_n_3236 = ~((mul_34_17_n_1737 & mul_34_17_n_2546) | (mul_34_17_n_2894 & mul_34_17_n_2522));
 assign mul_34_17_n_3235 = ((mul_34_17_n_1734 | mul_34_17_n_1918) & (mul_34_17_n_11588 | mul_34_17_n_1909));
 assign mul_34_17_n_3234 = ((mul_34_17_n_1736 | mul_34_17_n_2550) & (mul_34_17_n_11591 | mul_34_17_n_2554));
 assign mul_34_17_n_3232 = ~((mul_34_17_n_1751 & mul_34_17_n_2558) | (mul_34_17_n_2880 & mul_34_17_n_2580));
 assign mul_34_17_n_3231 = ~((mul_34_17_n_1741 & mul_34_17_n_1908) | (mul_34_17_n_2886 & mul_34_17_n_2700));
 assign mul_34_17_n_3230 = ~((mul_34_17_n_1745 & mul_34_17_n_2024) | (mul_34_17_n_2888 & mul_34_17_n_2185));
 assign mul_34_17_n_3228 = ~((mul_34_17_n_671 & mul_34_17_n_1067) | (mul_34_17_n_2918 & mul_34_17_n_1105));
 assign mul_34_17_n_3227 = ((mul_34_17_n_1740 | mul_34_17_n_1933) & (mul_34_17_n_11603 | mul_34_17_n_2030));
 assign mul_34_17_n_3226 = ((mul_34_17_n_1738 | mul_34_17_n_1910) & (mul_34_17_n_11606 | mul_34_17_n_1856));
 assign mul_34_17_n_3225 = ((mul_34_17_n_1746 | mul_34_17_n_2004) & (mul_34_17_n_11665 | mul_34_17_n_2227));
 assign mul_34_17_n_3224 = ((mul_34_17_n_1738 | mul_34_17_n_1854) & (mul_34_17_n_11606 | mul_34_17_n_2458));
 assign mul_34_17_n_3223 = ~((mul_34_17_n_681 & mul_34_17_n_839) | (mul_34_17_n_2928 & mul_34_17_n_843));
 assign mul_34_17_n_3222 = ~((mul_34_17_n_1753 & mul_34_17_n_1914) | (mul_34_17_n_2878 & mul_34_17_n_2524));
 assign mul_34_17_n_3221 = ((mul_34_17_n_1756 | mul_34_17_n_1576) & (mul_34_17_n_11582 | mul_34_17_n_866));
 assign mul_34_17_n_3220 = ~((mul_34_17_n_675 & mul_34_17_n_1001) | (mul_34_17_n_2922 & mul_34_17_n_975));
 assign mul_34_17_n_3219 = ((mul_34_17_n_678 | mul_34_17_n_894) & (mul_34_17_n_11543 | mul_34_17_n_891));
 assign mul_34_17_n_3218 = ~((mul_34_17_n_669 & mul_34_17_n_1157) | (mul_34_17_n_2916 & mul_34_17_n_1161));
 assign mul_34_17_n_3217 = ((mul_34_17_n_680 | mul_34_17_n_837) & (mul_34_17_n_11540 | mul_34_17_n_867));
 assign mul_34_17_n_3216 = ((mul_34_17_n_1756 | mul_34_17_n_1669) & (mul_34_17_n_11582 | mul_34_17_n_1770));
 assign mul_34_17_n_3215 = ~((mul_34_17_n_1742 | mul_34_17_n_2613) & (mul_34_17_n_11609 | mul_34_17_n_2566));
 assign mul_34_17_n_3214 = ((mul_34_17_n_1734 | mul_34_17_n_2607) & (mul_34_17_n_11588 | mul_34_17_n_1912));
 assign mul_34_17_n_3213 = ((mul_34_17_n_654 | mul_34_17_n_1625) & (mul_34_17_n_11579 | mul_34_17_n_1659));
 assign mul_34_17_n_3212 = ((mul_34_17_n_679 & mul_34_17_n_916) | (mul_34_17_n_2926 & mul_34_17_n_892));
 assign mul_34_17_n_3211 = ((mul_34_17_n_666 | mul_34_17_n_1188) & (mul_34_17_n_11561 | mul_34_17_n_1205));
 assign mul_34_17_n_3210 = ((mul_34_17_n_1736 | mul_34_17_n_1698) & (mul_34_17_n_11591 | mul_34_17_n_2207));
 assign mul_34_17_n_3209 = ((mul_34_17_n_1742 | mul_34_17_n_2634) & (mul_34_17_n_11609 | mul_34_17_n_2479));
 assign mul_34_17_n_3207 = ~((mul_34_17_n_1755 & mul_34_17_n_2477) | (mul_34_17_n_2898 & mul_34_17_n_2133));
 assign mul_34_17_n_3206 = ((mul_34_17_n_1750 | mul_34_17_n_2019) & (mul_34_17_n_11612 | mul_34_17_n_2582));
 assign mul_34_17_n_3205 = ~((mul_34_17_n_1737 & mul_34_17_n_2553) | (mul_34_17_n_2894 & mul_34_17_n_2222));
 assign mul_34_17_n_3204 = ((mul_34_17_n_658 | mul_34_17_n_1454) & (mul_34_17_n_11573 | mul_34_17_n_1485));
 assign mul_34_17_n_3202 = ((mul_34_17_n_1746 | mul_34_17_n_2087) & (mul_34_17_n_11678 | mul_34_17_n_2004));
 assign mul_34_17_n_3200 = ((mul_34_17_n_1740 | mul_34_17_n_1895) & (mul_34_17_n_11603 | mul_34_17_n_2048));
 assign mul_34_17_n_3198 = ~((mul_34_17_n_1751 & mul_34_17_n_2669) | (mul_34_17_n_2880 & mul_34_17_n_2599));
 assign mul_34_17_n_3197 = ((mul_34_17_n_682 | mul_34_17_n_826) & (mul_34_17_n_11537 | mul_34_17_n_829));
 assign mul_34_17_n_3195 = ((mul_34_17_n_672 | mul_34_17_n_1032) & (mul_34_17_n_11552 | mul_34_17_n_1035));
 assign mul_34_17_n_3194 = ~((mul_34_17_n_677 & mul_34_17_n_933) | (mul_34_17_n_2924 & mul_34_17_n_932));
 assign mul_34_17_n_3193 = ((mul_34_17_n_1748 | mul_34_17_n_2302) & (mul_34_17_n_11597 | mul_34_17_n_2132));
 assign mul_34_17_n_3192 = ~((mul_34_17_n_1751 & mul_34_17_n_2213) | (mul_34_17_n_2880 & mul_34_17_n_2584));
 assign mul_34_17_n_3191 = ((mul_34_17_n_1738 | mul_34_17_n_2685) & (mul_34_17_n_11606 | mul_34_17_n_1911));
 assign mul_34_17_n_3190 = ~((mul_34_17_n_1738 | mul_34_17_n_2098) & (mul_34_17_n_11606 | mul_34_17_n_1949));
 assign mul_34_17_n_3189 = ~((mul_34_17_n_667 & mul_34_17_n_1187) | (mul_34_17_n_2914 & mul_34_17_n_1218));
 assign mul_34_17_n_3188 = ((mul_34_17_n_1740 | mul_34_17_n_2144) & (mul_34_17_n_11603 | mul_34_17_n_1895));
 assign mul_34_17_n_3187 = ((mul_34_17_n_678 | mul_34_17_n_897) & (mul_34_17_n_11543 | mul_34_17_n_884));
 assign mul_34_17_n_3186 = ((mul_34_17_n_672 | mul_34_17_n_1056) & (mul_34_17_n_11552 | mul_34_17_n_1027));
 assign mul_34_17_n_3185 = ((mul_34_17_n_670 | mul_34_17_n_1068) & (mul_34_17_n_11555 | mul_34_17_n_1081));
 assign mul_34_17_n_3184 = ~((mul_34_17_n_675 & mul_34_17_n_979) | (mul_34_17_n_2922 & mul_34_17_n_986));
 assign mul_34_17_n_3183 = ~((mul_34_17_n_691 & mul_34_17_n_751) | (mul_34_17_n_2936 & mul_34_17_n_753));
 assign mul_34_17_n_3182 = ~((mul_34_17_n_1749 & mul_34_17_n_2337) | (mul_34_17_n_2890 & mul_34_17_n_1928));
 assign mul_34_17_n_3180 = ((mul_34_17_n_658 | mul_34_17_n_1488) & (mul_34_17_n_11573 | mul_34_17_n_1466));
 assign mul_34_17_n_3179 = ((mul_34_17_n_1746 | mul_34_17_n_1893) & (mul_34_17_n_11676 | mul_34_17_n_2087));
 assign mul_34_17_n_3178 = ((mul_34_17_n_1754 | mul_34_17_n_1881) & (mul_34_17_n_11585 | mul_34_17_n_2656));
 assign mul_34_17_n_3177 = ((mul_34_17_n_1750 | mul_34_17_n_2129) & (mul_34_17_n_11612 | mul_34_17_n_1954));
 assign mul_34_17_n_3176 = ~((mul_34_17_n_1757 & mul_34_17_n_799) | (mul_34_17_n_2900 & mul_34_17_n_2658));
 assign mul_34_17_n_3175 = ((mul_34_17_n_1734 | mul_34_17_n_2284) & (mul_34_17_n_11588 | mul_34_17_n_1922));
 assign mul_34_17_n_3174 = ((mul_34_17_n_1750 | mul_34_17_n_2032) & (mul_34_17_n_11612 | mul_34_17_n_2559));
 assign mul_34_17_n_3173 = ~((mul_34_17_n_657 & mul_34_17_n_1556) | (mul_34_17_n_2904 & mul_34_17_n_1574));
 assign mul_34_17_n_3172 = ~(mul_34_17_n_2856 ^ mul_34_17_n_2948);
 assign mul_34_17_n_3171 = ((mul_34_17_n_1738 | mul_34_17_n_2263) & (mul_34_17_n_11606 | mul_34_17_n_1996));
 assign mul_34_17_n_3170 = ((mul_34_17_n_656 | mul_34_17_n_1565) & (mul_34_17_n_11576 | mul_34_17_n_1536));
 assign mul_34_17_n_3169 = ~((mul_34_17_n_661 & mul_34_17_n_1397) | (mul_34_17_n_2908 & mul_34_17_n_1431));
 assign mul_34_17_n_3168 = ~((mul_34_17_n_656 | mul_34_17_n_1562) & (mul_34_17_n_11576 | mul_34_17_n_1542));
 assign mul_34_17_n_3166 = ((mul_34_17_n_1740 | mul_34_17_n_2660) & (mul_34_17_n_11603 | mul_34_17_n_2537));
 assign mul_34_17_n_3164 = ((mul_34_17_n_1746 | mul_34_17_n_2398) & (mul_34_17_n_11673 | mul_34_17_n_1893));
 assign mul_34_17_n_3162 = ((mul_34_17_n_1734 | mul_34_17_n_2150) & (mul_34_17_n_11588 | mul_34_17_n_2510));
 assign mul_34_17_n_3160 = ((mul_34_17_n_654 | mul_34_17_n_1651) & (mul_34_17_n_11579 | mul_34_17_n_1638));
 assign mul_34_17_n_3159 = ((mul_34_17_n_660 | mul_34_17_n_1412) & (mul_34_17_n_11570 | mul_34_17_n_1382));
 assign mul_34_17_n_3158 = ((mul_34_17_n_1738 | mul_34_17_n_2188) & (mul_34_17_n_11606 | mul_34_17_n_2110));
 assign mul_34_17_n_3157 = ((mul_34_17_n_662 | mul_34_17_n_1355) & (mul_34_17_n_11567 | mul_34_17_n_1368));
 assign mul_34_17_n_3156 = ((mul_34_17_n_1740 | mul_34_17_n_2699) & (mul_34_17_n_11603 | mul_34_17_n_2144));
 assign mul_34_17_n_3155 = ((mul_34_17_n_1736 | mul_34_17_n_2277) & (mul_34_17_n_11591 | mul_34_17_n_2346));
 assign mul_34_17_n_3154 = ((mul_34_17_n_1746 | mul_34_17_n_2335) & (mul_34_17_n_11675 | mul_34_17_n_2398));
 assign mul_34_17_n_3152 = ((mul_34_17_n_1750 | mul_34_17_n_1857) & (mul_34_17_n_11612 | mul_34_17_n_2089));
 assign mul_34_17_n_3151 = ((mul_34_17_n_1735 & mul_34_17_n_2074) | (mul_34_17_n_2896 & mul_34_17_n_2218));
 assign mul_34_17_n_3150 = ~((mul_34_17_n_1746 | mul_34_17_n_2412) & (mul_34_17_n_11680 | mul_34_17_n_2283));
 assign mul_34_17_n_3149 = ~((mul_34_17_n_659 & mul_34_17_n_1456) | (mul_34_17_n_2906 & mul_34_17_n_1512));
 assign mul_34_17_n_3148 = ((mul_34_17_n_1752 | mul_34_17_n_1983) & (mul_34_17_n_11615 | mul_34_17_n_2012));
 assign mul_34_17_n_3147 = ((mul_34_17_n_1756 | mul_34_17_n_1687) & (mul_34_17_n_11582 | mul_34_17_n_1677));
 assign mul_34_17_n_3145 = ((mul_34_17_n_1734 | mul_34_17_n_1997) & (mul_34_17_n_11588 | mul_34_17_n_1852));
 assign mul_34_17_n_3143 = ((mul_34_17_n_1734 | mul_34_17_n_1852) & (mul_34_17_n_11588 | mul_34_17_n_2150));
 assign mul_34_17_n_3141 = ~((mul_34_17_n_1737 & mul_34_17_n_2627) | (mul_34_17_n_2894 & mul_34_17_n_2464));
 assign mul_34_17_n_3140 = ~(mul_34_17_n_2946 ^ mul_34_17_n_2858);
 assign mul_34_17_n_3139 = ~((mul_34_17_n_675 & mul_34_17_n_977) | (mul_34_17_n_2922 & mul_34_17_n_969));
 assign mul_34_17_n_3137 = ((mul_34_17_n_1742 | mul_34_17_n_1879) & (mul_34_17_n_11609 | mul_34_17_n_2613));
 assign mul_34_17_n_3135 = ((mul_34_17_n_1756 | mul_34_17_n_1667) & (mul_34_17_n_11582 | mul_34_17_n_1974));
 assign mul_34_17_n_3134 = ((mul_34_17_n_1742 | mul_34_17_n_2166) & (mul_34_17_n_11609 | mul_34_17_n_2229));
 assign mul_34_17_n_3132 = ~((mul_34_17_n_1743 & mul_34_17_n_2238) | (mul_34_17_n_2882 & mul_34_17_n_2275));
 assign mul_34_17_n_3130 = ((mul_34_17_n_1740 | mul_34_17_n_1913) & (mul_34_17_n_11603 | mul_34_17_n_2079));
 assign mul_34_17_n_3128 = ((mul_34_17_n_1748 | mul_34_17_n_1861) & (mul_34_17_n_11597 | mul_34_17_n_2549));
 assign mul_34_17_n_3127 = ((mul_34_17_n_658 | mul_34_17_n_1515) & (mul_34_17_n_11573 | mul_34_17_n_1463));
 assign mul_34_17_n_3126 = ((mul_34_17_n_1754 | mul_34_17_n_2548) & (mul_34_17_n_11585 | mul_34_17_n_1916));
 assign mul_34_17_n_3125 = ~((mul_34_17_n_1743 & mul_34_17_n_2609) | (mul_34_17_n_2882 & mul_34_17_n_2612));
 assign mul_34_17_n_3124 = ((mul_34_17_n_684 | mul_34_17_n_797) & (mul_34_17_n_11534 | mul_34_17_n_786));
 assign mul_34_17_n_3123 = ((mul_34_17_n_1748 | mul_34_17_n_2132) & (mul_34_17_n_11597 | mul_34_17_n_2357));
 assign mul_34_17_n_3122 = ((mul_34_17_n_664 | mul_34_17_n_1295) & (mul_34_17_n_11564 | mul_34_17_n_1276));
 assign mul_34_17_n_3121 = ~((mul_34_17_n_685 & mul_34_17_n_794) | (mul_34_17_n_2931 & mul_34_17_n_779));
 assign mul_34_17_n_3120 = ((mul_34_17_n_664 | mul_34_17_n_1271) & (mul_34_17_n_11564 | mul_34_17_n_1278));
 assign mul_34_17_n_3119 = ~((mul_34_17_n_657 & mul_34_17_n_1564) | (mul_34_17_n_2904 & mul_34_17_n_1521));
 assign mul_34_17_n_3118 = ~(mul_34_17_n_3001 | mul_34_17_n_2748);
 assign mul_34_17_n_3117 = ((mul_34_17_n_1750 | mul_34_17_n_1855) & (mul_34_17_n_11612 | mul_34_17_n_2500));
 assign mul_34_17_n_3115 = ~((mul_34_17_n_680 | mul_34_17_n_846) & (mul_34_17_n_11540 | mul_34_17_n_857));
 assign mul_34_17_n_3113 = ~((mul_34_17_n_679 & mul_34_17_n_909) | (mul_34_17_n_2926 & mul_34_17_n_915));
 assign mul_34_17_n_3112 = ((mul_34_17_n_1756 | mul_34_17_n_1476) & (mul_34_17_n_11582 | mul_34_17_n_903));
 assign mul_34_17_n_3111 = ((mul_34_17_n_1752 | mul_34_17_n_2353) & (mul_34_17_n_11615 | mul_34_17_n_2136));
 assign mul_34_17_n_3109 = ~((mul_34_17_n_1757 & mul_34_17_n_1765) | (mul_34_17_n_2900 & mul_34_17_n_1626));
 assign mul_34_17_n_3108 = ((mul_34_17_n_676 | mul_34_17_n_959) & (mul_34_17_n_11546 | mul_34_17_n_941));
 assign mul_34_17_n_3107 = ((mul_34_17_n_680 | mul_34_17_n_847) & (mul_34_17_n_11540 | mul_34_17_n_849));
 assign mul_34_17_n_3106 = ~((mul_34_17_n_691 & mul_34_17_n_746) | (mul_34_17_n_2936 & mul_34_17_n_710));
 assign mul_34_17_n_3105 = ((mul_34_17_n_666 | mul_34_17_n_1209) & (mul_34_17_n_11561 | mul_34_17_n_1211));
 assign mul_34_17_n_3104 = ~((mul_34_17_n_1739 & mul_34_17_n_1847) | (mul_34_17_n_2884 & mul_34_17_n_2126));
 assign mul_34_17_n_3103 = ~((mul_34_17_n_1741 & mul_34_17_n_2157) | (mul_34_17_n_2886 & mul_34_17_n_2193));
 assign mul_34_17_n_3102 = ~((mul_34_17_n_1745 & mul_34_17_n_1691) | (mul_34_17_n_2888 & mul_34_17_n_2463));
 assign mul_34_17_n_3101 = ((mul_34_17_n_659 & mul_34_17_n_1506) | (mul_34_17_n_2906 & mul_34_17_n_1448));
 assign mul_34_17_n_3099 = ((mul_34_17_n_660 | mul_34_17_n_1378) & (mul_34_17_n_11570 | mul_34_17_n_1443));
 assign mul_34_17_n_3098 = ((mul_34_17_n_1734 | mul_34_17_n_2516) & (mul_34_17_n_11588 | mul_34_17_n_1892));
 assign mul_34_17_n_3097 = ((mul_34_17_n_1755 & mul_34_17_n_1849) | (mul_34_17_n_2898 & mul_34_17_n_2252));
 assign mul_34_17_n_3096 = ((mul_34_17_n_680 | mul_34_17_n_864) & (mul_34_17_n_11540 | mul_34_17_n_837));
 assign mul_34_17_n_3094 = ((mul_34_17_n_682 | mul_34_17_n_801) & (mul_34_17_n_11537 | mul_34_17_n_811));
 assign mul_34_17_n_3093 = ~((mul_34_17_n_1753 & mul_34_17_n_2306) | (mul_34_17_n_2878 & mul_34_17_n_2338));
 assign mul_34_17_n_3092 = ((mul_34_17_n_1748 | mul_34_17_n_2294) & (mul_34_17_n_11597 | mul_34_17_n_2076));
 assign mul_34_17_n_3091 = ((mul_34_17_n_1752 | mul_34_17_n_2400) & (mul_34_17_n_11615 | mul_34_17_n_2172));
 assign mul_34_17_n_3089 = ~((mul_34_17_n_675 & mul_34_17_n_973) | (mul_34_17_n_2922 & mul_34_17_n_988));
 assign mul_34_17_n_3088 = ((mul_34_17_n_680 | mul_34_17_n_834) & (mul_34_17_n_11540 | mul_34_17_n_846));
 assign mul_34_17_n_3087 = ((mul_34_17_n_1745 & mul_34_17_n_2482) | (mul_34_17_n_2888 & mul_34_17_n_2689));
 assign mul_34_17_n_3086 = ~((mul_34_17_n_687 & mul_34_17_n_695) | (mul_34_17_n_2933 & mul_34_17_n_739));
 assign mul_34_17_n_3085 = ((mul_34_17_n_1756 | mul_34_17_n_1665) & (mul_34_17_n_11582 | mul_34_17_n_1684));
 assign mul_34_17_n_3084 = ((mul_34_17_n_1754 | mul_34_17_n_1844) & (mul_34_17_n_11585 | mul_34_17_n_1842));
 assign mul_34_17_n_3083 = ((mul_34_17_n_1748 | mul_34_17_n_2556) & (mul_34_17_n_11597 | mul_34_17_n_2230));
 assign mul_34_17_n_3082 = ((mul_34_17_n_1747 & mul_34_17_n_1936) | (mul_34_17_n_11593 & mul_34_17_n_2108));
 assign mul_34_17_n_3080 = ((mul_34_17_n_656 | mul_34_17_n_1568) & (mul_34_17_n_11576 | mul_34_17_n_1546));
 assign mul_34_17_n_3079 = ((mul_34_17_n_682 | mul_34_17_n_802) & (mul_34_17_n_11537 | mul_34_17_n_1701));
 assign mul_34_17_n_3078 = ((mul_34_17_n_1734 | mul_34_17_n_2171) & (mul_34_17_n_11588 | mul_34_17_n_2520));
 assign mul_34_17_n_3076 = ((mul_34_17_n_662 | mul_34_17_n_1373) & (mul_34_17_n_11567 | mul_34_17_n_1361));
 assign mul_34_17_n_3075 = ((mul_34_17_n_1751 & mul_34_17_n_2134) | (mul_34_17_n_2880 & mul_34_17_n_1960));
 assign mul_34_17_n_3074 = ((mul_34_17_n_662 | mul_34_17_n_1353) & (mul_34_17_n_11567 | mul_34_17_n_1356));
 assign mul_34_17_n_3072 = ~((mul_34_17_n_674 | mul_34_17_n_982) & (mul_34_17_n_11549 | mul_34_17_n_987));
 assign mul_34_17_n_3070 = ~((mul_34_17_n_687 & mul_34_17_n_747) | (mul_34_17_n_2933 & mul_34_17_n_807));
 assign mul_34_17_n_3069 = ((mul_34_17_n_670 | mul_34_17_n_1081) & (mul_34_17_n_11555 | mul_34_17_n_1097));
 assign mul_34_17_n_3068 = ~((mul_34_17_n_685 & mul_34_17_n_777) | (mul_34_17_n_2931 & mul_34_17_n_795));
 assign mul_34_17_n_3065 = ~((mul_34_17_n_1753 & mul_34_17_n_2359) | (mul_34_17_n_2878 & mul_34_17_n_2023));
 assign mul_34_17_n_3063 = ((mul_34_17_n_1742 | mul_34_17_n_2496) & (mul_34_17_n_11609 | mul_34_17_n_2214));
 assign mul_34_17_n_3062 = ~((mul_34_17_n_654 | mul_34_17_n_1629) & (mul_34_17_n_11579 | mul_34_17_n_1631));
 assign mul_34_17_n_3061 = ((mul_34_17_n_664 | mul_34_17_n_1284) & (mul_34_17_n_11564 | mul_34_17_n_1296));
 assign mul_34_17_n_3059 = ~(mul_34_17_n_2861 ^ mul_34_17_n_2943);
 assign mul_34_17_n_3058 = ~((mul_34_17_n_675 & mul_34_17_n_968) | (mul_34_17_n_2922 & mul_34_17_n_990));
 assign mul_34_17_n_3057 = ((mul_34_17_n_1749 & mul_34_17_n_2684) | (mul_34_17_n_2890 & mul_34_17_n_2122));
 assign mul_34_17_n_3056 = ~((mul_34_17_n_1744 | mul_34_17_n_2399) & (mul_34_17_n_11600 | mul_34_17_n_2073));
 assign mul_34_17_n_3055 = ((mul_34_17_n_668 | mul_34_17_n_1146) & (mul_34_17_n_11558 | mul_34_17_n_1128));
 assign mul_34_17_n_3054 = ~((mul_34_17_n_1734 | mul_34_17_n_2031) & (mul_34_17_n_11588 | mul_34_17_n_1941));
 assign mul_34_17_n_3053 = ~((mul_34_17_n_666 | mul_34_17_n_1207) & (mul_34_17_n_11561 | mul_34_17_n_1213));
 assign mul_34_17_n_3038 = ~mul_34_17_n_3039;
 assign mul_34_17_n_3035 = ~mul_34_17_n_3034;
 assign mul_34_17_n_3025 = ~mul_34_17_n_3026;
 assign mul_34_17_n_3024 = ~mul_34_17_n_3006;
 assign mul_34_17_n_3021 = ~(mul_34_17_n_11552 | mul_34_17_n_469);
 assign mul_34_17_n_3020 = ~(mul_34_17_n_11570 | mul_34_17_n_456);
 assign mul_34_17_n_3019 = ~(mul_34_17_n_11567 | mul_34_17_n_458);
 assign mul_34_17_n_3018 = ~(mul_34_17_n_11564 | mul_34_17_n_461);
 assign mul_34_17_n_3017 = ~(mul_34_17_n_11561 | mul_34_17_n_463);
 assign mul_34_17_n_3016 = ~(mul_34_17_n_11558 | mul_34_17_n_464);
 assign mul_34_17_n_3015 = ~(mul_34_17_n_11555 | mul_34_17_n_467);
 assign mul_34_17_n_3014 = ~(mul_34_17_n_11573 | mul_34_17_n_453);
 assign mul_34_17_n_3013 = ~(mul_34_17_n_11549 | mul_34_17_n_471);
 assign mul_34_17_n_3012 = ~(mul_34_17_n_11546 | mul_34_17_n_472);
 assign mul_34_17_n_3011 = ~(mul_34_17_n_11543 | mul_34_17_n_475);
 assign mul_34_17_n_3010 = ~(mul_34_17_n_11540 | mul_34_17_n_477);
 assign mul_34_17_n_3009 = ~(mul_34_17_n_11534 | mul_34_17_n_479);
 assign mul_34_17_n_3008 = ~(mul_34_17_n_11531 | mul_34_17_n_482);
 assign mul_34_17_n_3007 = ~(mul_34_17_n_11525 | mul_34_17_n_484);
 assign mul_34_17_n_3041 = ~(mul_34_17_n_2859 | mul_34_17_n_2947);
 assign mul_34_17_n_3040 = ~(mul_34_17_n_2862 | mul_34_17_n_2943);
 assign mul_34_17_n_3039 = ~(mul_34_17_n_2871 | mul_34_17_n_2239);
 assign mul_34_17_n_3037 = ~(mul_34_17_n_2850 | mul_34_17_n_2938);
 assign mul_34_17_n_3036 = ~(mul_34_17_n_2863 | mul_34_17_n_2941);
 assign mul_34_17_n_3034 = ~(mul_34_17_n_2860 | mul_34_17_n_2949);
 assign mul_34_17_n_3033 = ~(mul_34_17_n_2857 | mul_34_17_n_2948);
 assign mul_34_17_n_3032 = ~(mul_34_17_n_2874 | mul_34_17_n_2950);
 assign mul_34_17_n_3031 = ~(mul_34_17_n_2858 | mul_34_17_n_2946);
 assign mul_34_17_n_3030 = ~(mul_34_17_n_2869 | mul_34_17_n_2955);
 assign mul_34_17_n_3029 = ~(mul_34_17_n_2870 | mul_34_17_n_2952);
 assign mul_34_17_n_3028 = ~(mul_34_17_n_2864 | mul_34_17_n_2969);
 assign mul_34_17_n_3027 = ~(mul_34_17_n_2866 | mul_34_17_n_2956);
 assign mul_34_17_n_3026 = ~(mul_34_17_n_2829 | mul_34_17_n_2940);
 assign mul_34_17_n_3006 = ~(mul_34_17_n_2875 | mul_34_17_n_2966);
 assign mul_34_17_n_3023 = ~(mul_34_17_n_2877 | mul_34_17_n_2964);
 assign mul_34_17_n_3022 = ~(mul_34_17_n_2873 | mul_34_17_n_2967);
 assign mul_34_17_n_3005 = ~mul_34_17_n_2978;
 assign mul_34_17_n_2994 = ~mul_34_17_n_2974;
 assign mul_34_17_n_2992 = ~mul_34_17_n_2972;
 assign mul_34_17_n_2990 = ~(mul_34_17_n_11582 | mul_34_17_n_447);
 assign mul_34_17_n_2989 = ~(mul_34_17_n_11597 | mul_34_17_n_442);
 assign mul_34_17_n_2988 = ~(mul_34_17_n_11600 | mul_34_17_n_446);
 assign mul_34_17_n_2987 = ~(mul_34_17_n_11609 | mul_34_17_n_429);
 assign mul_34_17_n_2986 = ~(mul_34_17_n_11588 | mul_34_17_n_443);
 assign mul_34_17_n_2985 = ~(mul_34_17_n_11615 | mul_34_17_n_439);
 assign mul_34_17_n_2984 = ~(mul_34_17_n_11694 | mul_34_17_n_427);
 assign mul_34_17_n_2983 = ~(mul_34_17_n_11612 | mul_34_17_n_440);
 assign mul_34_17_n_2982 = ~(mul_34_17_n_11603 | mul_34_17_n_438);
 assign mul_34_17_n_2981 = ~(mul_34_17_n_11606 | mul_34_17_n_441);
 assign mul_34_17_n_2980 = ~(mul_34_17_n_11591 | mul_34_17_n_431);
 assign mul_34_17_n_2979 = ~(mul_34_17_n_11585 | mul_34_17_n_455);
 assign mul_34_17_n_2978 = ~(mul_34_17_n_2846 | mul_34_17_n_2720);
 assign mul_34_17_n_2977 = ~(mul_34_17_n_11576 | mul_34_17_n_451);
 assign mul_34_17_n_3004 = ~(mul_34_17_n_2846 & mul_34_17_n_2720);
 assign mul_34_17_n_3003 = ~(mul_34_17_n_11540 | mul_34_17_n_868);
 assign mul_34_17_n_3002 = ~(mul_34_17_n_11561 | mul_34_17_n_1241);
 assign mul_34_17_n_3001 = ~(mul_34_17_n_11558 | mul_34_17_n_1137);
 assign mul_34_17_n_3000 = ~(mul_34_17_n_11558 | mul_34_17_n_1140);
 assign mul_34_17_n_2976 = ~(mul_34_17_n_2904 & mul_34_17_n_1573);
 assign mul_34_17_n_2999 = ~(mul_34_17_n_11573 | mul_34_17_n_1486);
 assign mul_34_17_n_2998 = ~(mul_34_17_n_11612 | mul_34_17_n_2325);
 assign mul_34_17_n_2975 = ~(mul_34_17_n_2922 & mul_34_17_n_1012);
 assign mul_34_17_n_2997 = ~(mul_34_17_n_11579 | mul_34_17_n_1629);
 assign mul_34_17_n_2996 = ~(mul_34_17_n_11591 | mul_34_17_n_1896);
 assign mul_34_17_n_2995 = ~(mul_34_17_n_2906 & mul_34_17_n_1495);
 assign mul_34_17_n_2974 = ~(mul_34_17_n_11528 | mul_34_17_n_706);
 assign mul_34_17_n_2993 = ~(mul_34_17_n_11600 | mul_34_17_n_2637);
 assign mul_34_17_n_2973 = ~(mul_34_17_n_11579 | mul_34_17_n_450);
 assign mul_34_17_n_2972 = ~(mul_34_17_n_2868 & mul_34_17_n_2743);
 assign mul_34_17_n_2970 = ~(mul_34_17_n_2868 | mul_34_17_n_2743);
 assign mul_34_17_n_2945 = ~mul_34_17_n_2944;
 assign mul_34_17_n_2936 = ~mul_34_17_n_11525;
 assign mul_34_17_n_2933 = ~mul_34_17_n_11531;
 assign mul_34_17_n_2931 = ~mul_34_17_n_11534;
 assign mul_34_17_n_2928 = ~mul_34_17_n_11540;
 assign mul_34_17_n_2926 = ~mul_34_17_n_11543;
 assign mul_34_17_n_2924 = ~mul_34_17_n_11546;
 assign mul_34_17_n_2922 = ~mul_34_17_n_11549;
 assign mul_34_17_n_2920 = ~mul_34_17_n_11552;
 assign mul_34_17_n_2918 = ~mul_34_17_n_11555;
 assign mul_34_17_n_2916 = ~mul_34_17_n_11558;
 assign mul_34_17_n_2914 = ~mul_34_17_n_11561;
 assign mul_34_17_n_2912 = ~mul_34_17_n_11564;
 assign mul_34_17_n_2910 = ~mul_34_17_n_11567;
 assign mul_34_17_n_2908 = ~mul_34_17_n_11570;
 assign mul_34_17_n_2906 = ~mul_34_17_n_11573;
 assign mul_34_17_n_2904 = ~mul_34_17_n_11576;
 assign mul_34_17_n_2902 = ~mul_34_17_n_11579;
 assign mul_34_17_n_2900 = ~mul_34_17_n_11582;
 assign mul_34_17_n_2898 = ~mul_34_17_n_11585;
 assign mul_34_17_n_2896 = ~mul_34_17_n_11588;
 assign mul_34_17_n_2894 = ~mul_34_17_n_11591;
 assign mul_34_17_n_2890 = ~mul_34_17_n_11597;
 assign mul_34_17_n_2888 = ~mul_34_17_n_11600;
 assign mul_34_17_n_2886 = ~mul_34_17_n_11603;
 assign mul_34_17_n_2884 = ~mul_34_17_n_11606;
 assign mul_34_17_n_2882 = ~mul_34_17_n_11609;
 assign mul_34_17_n_2880 = ~mul_34_17_n_11612;
 assign mul_34_17_n_2878 = ~mul_34_17_n_11615;
 assign mul_34_17_n_2969 = ~(mul_34_17_n_2772 & mul_34_17_n_563);
 assign mul_34_17_n_2968 = ~(mul_34_17_n_2768 & mul_34_17_n_558);
 assign mul_34_17_n_2967 = ~(mul_34_17_n_2771 & mul_34_17_n_561);
 assign mul_34_17_n_2966 = ~(mul_34_17_n_2706 & mul_34_17_n_499);
 assign mul_34_17_n_2965 = ~(mul_34_17_n_2710 & mul_34_17_n_569);
 assign mul_34_17_n_2964 = ~(mul_34_17_n_2773 & mul_34_17_n_498);
 assign mul_34_17_n_2963 = ~(mul_34_17_n_2775 & mul_34_17_n_537);
 assign mul_34_17_n_2962 = ~(mul_34_17_n_2770 & mul_34_17_n_506);
 assign mul_34_17_n_2961 = ~(mul_34_17_n_2711 & mul_34_17_n_550);
 assign mul_34_17_n_2960 = ~(mul_34_17_n_2776 & mul_34_17_n_503);
 assign mul_34_17_n_2959 = ~(mul_34_17_n_2705 & mul_34_17_n_545);
 assign mul_34_17_n_2958 = ~(mul_34_17_n_2767 & mul_34_17_n_534);
 assign mul_34_17_n_2957 = ~(mul_34_17_n_2765 & mul_34_17_n_565);
 assign mul_34_17_n_2956 = ~(mul_34_17_n_2764 & mul_34_17_n_541);
 assign mul_34_17_n_2955 = ~(mul_34_17_n_2763 & mul_34_17_n_505);
 assign mul_34_17_n_2954 = ~(mul_34_17_n_2704 & mul_34_17_n_533);
 assign mul_34_17_n_2953 = ~(mul_34_17_n_2755 & mul_34_17_n_502);
 assign mul_34_17_n_2952 = ~(mul_34_17_n_2760 & mul_34_17_n_500);
 assign mul_34_17_n_2951 = ~(mul_34_17_n_2756 & mul_34_17_n_543);
 assign mul_34_17_n_2950 = ~(mul_34_17_n_2757 & mul_34_17_n_507);
 assign mul_34_17_n_2949 = ~(mul_34_17_n_2774 & mul_34_17_n_501);
 assign mul_34_17_n_2948 = ~(mul_34_17_n_2759 & mul_34_17_n_535);
 assign mul_34_17_n_2947 = ~(mul_34_17_n_2761 & mul_34_17_n_554);
 assign mul_34_17_n_2946 = ~(mul_34_17_n_2762 & mul_34_17_n_539);
 assign mul_34_17_n_2944 = ~(mul_34_17_n_2766 & mul_34_17_n_557);
 assign mul_34_17_n_2943 = ~(mul_34_17_n_2769 & mul_34_17_n_510);
 assign mul_34_17_n_2942 = ~(mul_34_17_n_2709 & mul_34_17_n_570);
 assign mul_34_17_n_2941 = ~(mul_34_17_n_2707 & mul_34_17_n_546);
 assign mul_34_17_n_2940 = ~(mul_34_17_n_2777 & mul_34_17_n_514);
 assign mul_34_17_n_2939 = ~(mul_34_17_n_2708 & mul_34_17_n_556);
 assign mul_34_17_n_2938 = ~(mul_34_17_n_2758 & mul_34_17_n_553);
 assign mul_34_17_n_2877 = ~mul_34_17_n_2876;
 assign mul_34_17_n_2872 = ~mul_34_17_n_2871;
 assign mul_34_17_n_2866 = ~mul_34_17_n_2865;
 assign mul_34_17_n_2862 = ~mul_34_17_n_2861;
 assign mul_34_17_n_2857 = ~mul_34_17_n_2856;
 assign mul_34_17_n_2810 = ~mul_34_17_n_2809;
 assign mul_34_17_n_2876 = ((mul_34_17_n_1809 & {in2[0]}) | (mul_34_17_n_1800 & mul_34_17_n_516));
 assign mul_34_17_n_2875 = ~((mul_34_17_n_1688 & {in2[0]}) | (mul_34_17_n_1795 & mul_34_17_n_516));
 assign mul_34_17_n_2874 = ~((mul_34_17_n_1838 & {in2[0]}) | (mul_34_17_n_1827 & mul_34_17_n_516));
 assign mul_34_17_n_2873 = ~((mul_34_17_n_1798 & {in2[0]}) | (mul_34_17_n_1796 & mul_34_17_n_516));
 assign mul_34_17_n_2871 = ~((mul_34_17_n_1824 & {in2[0]}) | (mul_34_17_n_1703 & mul_34_17_n_516));
 assign mul_34_17_n_2870 = ~((mul_34_17_n_1797 & {in2[0]}) | (mul_34_17_n_1813 & mul_34_17_n_516));
 assign mul_34_17_n_2869 = ~((mul_34_17_n_1802 & {in2[0]}) | (mul_34_17_n_1821 & mul_34_17_n_516));
 assign mul_34_17_n_2868 = ((mul_34_17_n_1810 & {in2[0]}) | (mul_34_17_n_1824 & mul_34_17_n_516));
 assign mul_34_17_n_2867 = ((mul_34_17_n_1784 & {in2[0]}) | (mul_34_17_n_1810 & mul_34_17_n_516));
 assign mul_34_17_n_2865 = ((mul_34_17_n_1825 & {in2[0]}) | (mul_34_17_n_1811 & mul_34_17_n_516));
 assign mul_34_17_n_2864 = ~((mul_34_17_n_1803 & {in2[0]}) | (mul_34_17_n_1805 & mul_34_17_n_516));
 assign mul_34_17_n_2863 = ~((mul_34_17_n_1789 & {in2[0]}) | (mul_34_17_n_1791 & mul_34_17_n_516));
 assign mul_34_17_n_2861 = ((mul_34_17_n_1804 & {in2[0]}) | (mul_34_17_n_1801 & mul_34_17_n_516));
 assign mul_34_17_n_2860 = ~((mul_34_17_n_1817 & {in2[0]}) | (mul_34_17_n_1793 & mul_34_17_n_516));
 assign mul_34_17_n_2859 = ~((mul_34_17_n_1794 & {in2[0]}) | (mul_34_17_n_1830 & mul_34_17_n_516));
 assign mul_34_17_n_2858 = ~((mul_34_17_n_1779 & {in2[0]}) | (mul_34_17_n_1785 & mul_34_17_n_516));
 assign mul_34_17_n_2856 = ((mul_34_17_n_1788 & {in2[0]}) | (mul_34_17_n_1834 & mul_34_17_n_516));
 assign mul_34_17_n_2855 = ~((mul_34_17_n_1793 & {in2[0]}) | (mul_34_17_n_1839 & mul_34_17_n_516));
 assign mul_34_17_n_2854 = ~((mul_34_17_n_1836 & {in2[0]}) | (mul_34_17_n_1838 & mul_34_17_n_516));
 assign mul_34_17_n_2853 = ~((mul_34_17_n_1778 & {in2[0]}) | (mul_34_17_n_1777 & mul_34_17_n_516));
 assign mul_34_17_n_2852 = ~((mul_34_17_n_1826 & {in2[0]}) | (mul_34_17_n_1822 & mul_34_17_n_516));
 assign mul_34_17_n_2851 = ~((mul_34_17_n_1805 & {in2[0]}) | (mul_34_17_n_1835 & mul_34_17_n_516));
 assign mul_34_17_n_2850 = ~((mul_34_17_n_1792 & {in2[0]}) | (mul_34_17_n_1829 & mul_34_17_n_516));
 assign mul_34_17_n_2849 = ((mul_34_17_n_1786 & {in2[0]}) | (mul_34_17_n_1836 & mul_34_17_n_516));
 assign mul_34_17_n_2848 = ~((mul_34_17_n_1807 & {in2[0]}) | (mul_34_17_n_1798 & mul_34_17_n_516));
 assign mul_34_17_n_2847 = ((mul_34_17_n_1816 & {in2[0]}) | (mul_34_17_n_1826 & mul_34_17_n_516));
 assign mul_34_17_n_2846 = ~((mul_34_17_n_1819 & {in2[0]}) | (mul_34_17_n_1784 & mul_34_17_n_516));
 assign mul_34_17_n_2845 = ~((mul_34_17_n_1785 & {in2[0]}) | (mul_34_17_n_1802 & mul_34_17_n_516));
 assign mul_34_17_n_2844 = ((mul_34_17_n_1800 & {in2[0]}) | (mul_34_17_n_1803 & mul_34_17_n_516));
 assign mul_34_17_n_2843 = ((mul_34_17_n_1780 & {in2[0]}) | (mul_34_17_n_1799 & mul_34_17_n_516));
 assign mul_34_17_n_2842 = ~((mul_34_17_n_1814 & {in2[0]}) | (mul_34_17_n_1778 & mul_34_17_n_516));
 assign mul_34_17_n_2841 = ~((mul_34_17_n_1801 & {in2[0]}) | (mul_34_17_n_1809 & mul_34_17_n_516));
 assign mul_34_17_n_2840 = ~((mul_34_17_n_1777 & {in2[0]}) | (mul_34_17_n_1790 & mul_34_17_n_516));
 assign mul_34_17_n_2839 = ~((mul_34_17_n_1830 & {in2[0]}) | (mul_34_17_n_1779 & mul_34_17_n_516));
 assign mul_34_17_n_2838 = ~((mul_34_17_n_1799 & {in2[0]}) | (mul_34_17_n_1783 & mul_34_17_n_516));
 assign mul_34_17_n_2837 = ((mul_34_17_n_1790 & {in2[0]}) | (mul_34_17_n_1787 & mul_34_17_n_516));
 assign mul_34_17_n_2836 = ((mul_34_17_n_1822 & {in2[0]}) | (mul_34_17_n_1806 & mul_34_17_n_516));
 assign mul_34_17_n_2835 = ~((mul_34_17_n_1781 & {in2[0]}) | (mul_34_17_n_1782 & mul_34_17_n_516));
 assign mul_34_17_n_2834 = ~((mul_34_17_n_1808 & {in2[0]}) | (mul_34_17_n_1815 & mul_34_17_n_516));
 assign mul_34_17_n_2833 = ~((mul_34_17_n_1815 & {in2[0]}) | (mul_34_17_n_1817 & mul_34_17_n_516));
 assign mul_34_17_n_2832 = ~((mul_34_17_n_1821 & {in2[0]}) | (mul_34_17_n_1825 & mul_34_17_n_516));
 assign mul_34_17_n_2831 = ~((mul_34_17_n_1834 & {in2[0]}) | (mul_34_17_n_1797 & mul_34_17_n_516));
 assign mul_34_17_n_2830 = ~((mul_34_17_n_1812 & {in2[0]}) | (mul_34_17_n_1786 & mul_34_17_n_516));
 assign mul_34_17_n_2829 = ~((mul_34_17_n_1839 & {in2[0]}) | (mul_34_17_n_1819 & mul_34_17_n_516));
 assign mul_34_17_n_2828 = ~((mul_34_17_n_1837 & {in2[0]}) | (mul_34_17_n_1808 & mul_34_17_n_516));
 assign mul_34_17_n_2827 = ((mul_34_17_n_1782 & {in2[0]}) | (mul_34_17_n_1807 & mul_34_17_n_516));
 assign mul_34_17_n_2826 = ~((mul_34_17_n_1806 & {in2[0]}) | (mul_34_17_n_1780 & mul_34_17_n_516));
 assign mul_34_17_n_2825 = ~((mul_34_17_n_1811 & {in2[0]}) | (mul_34_17_n_1818 & mul_34_17_n_516));
 assign mul_34_17_n_2824 = ~((mul_34_17_n_1795 & {in2[0]}) | (mul_34_17_n_1789 & mul_34_17_n_516));
 assign mul_34_17_n_2823 = ~((mul_34_17_n_1818 & {in2[0]}) | (mul_34_17_n_1820 & mul_34_17_n_516));
 assign mul_34_17_n_2822 = ~((mul_34_17_n_1813 & {in2[0]}) | (mul_34_17_n_1794 & mul_34_17_n_516));
 assign mul_34_17_n_2821 = ~((mul_34_17_n_1796 & {in2[0]}) | (mul_34_17_n_1804 & mul_34_17_n_516));
 assign mul_34_17_n_2820 = ((mul_34_17_n_1835 & {in2[0]}) | (mul_34_17_n_1837 & mul_34_17_n_516));
 assign mul_34_17_n_2819 = ~((mul_34_17_n_1783 & {in2[0]}) | (mul_34_17_n_1812 & mul_34_17_n_516));
 assign mul_34_17_n_2818 = ~((mul_34_17_n_1787 & {in2[0]}) | (mul_34_17_n_1823 & mul_34_17_n_516));
 assign mul_34_17_n_2817 = ~((mul_34_17_n_1820 & {in2[0]}) | (mul_34_17_n_1828 & mul_34_17_n_516));
 assign mul_34_17_n_2816 = ((mul_34_17_n_1832 & {in2[0]}) | (mul_34_17_n_1781 & mul_34_17_n_516));
 assign mul_34_17_n_2815 = ~((mul_34_17_n_1833 & {in2[0]}) | (mul_34_17_n_1832 & mul_34_17_n_516));
 assign mul_34_17_n_2814 = ~((mul_34_17_n_1827 & {in2[0]}) | (mul_34_17_n_1792 & mul_34_17_n_516));
 assign mul_34_17_n_2813 = ((mul_34_17_n_1828 & {in2[0]}) | (mul_34_17_n_1833 & mul_34_17_n_516));
 assign mul_34_17_n_2812 = ~((mul_34_17_n_1829 & {in2[0]}) | (mul_34_17_n_1788 & mul_34_17_n_516));
 assign mul_34_17_n_2811 = ~((mul_34_17_n_1823 & {in2[0]}) | (mul_34_17_n_1816 & mul_34_17_n_516));
 assign mul_34_17_n_2809 = ((mul_34_17_n_1791 & {in2[0]}) | (mul_34_17_n_1814 & mul_34_17_n_516));
 assign mul_34_17_n_2777 = ~(mul_34_17_n_1715 | mul_34_17_n_412);
 assign mul_34_17_n_2776 = ~(mul_34_17_n_1711 | mul_34_17_n_417);
 assign mul_34_17_n_2775 = ~(mul_34_17_n_1725 | mul_34_17_n_418);
 assign mul_34_17_n_2774 = ~(mul_34_17_n_1717 | mul_34_17_n_396);
 assign mul_34_17_n_2773 = ~(mul_34_17_n_1719 | mul_34_17_n_393);
 assign mul_34_17_n_2772 = ~(mul_34_17_n_1729 | mul_34_17_n_394);
 assign mul_34_17_n_2771 = ~(mul_34_17_n_1706 | mul_34_17_n_395);
 assign mul_34_17_n_2770 = ~(mul_34_17_n_1724 | mul_34_17_n_416);
 assign mul_34_17_n_2769 = ~(mul_34_17_n_1716 | mul_34_17_n_415);
 assign mul_34_17_n_2768 = ~(mul_34_17_n_1730 | mul_34_17_n_414);
 assign mul_34_17_n_2767 = ~(mul_34_17_n_1733 | mul_34_17_n_398);
 assign mul_34_17_n_2766 = ~(mul_34_17_n_1718 | mul_34_17_n_413);
 assign mul_34_17_n_2765 = ~(mul_34_17_n_1723 | mul_34_17_n_399);
 assign mul_34_17_n_2764 = ~(mul_34_17_n_1721 | mul_34_17_n_400);
 assign mul_34_17_n_2763 = ~(mul_34_17_n_1710 | mul_34_17_n_401);
 assign mul_34_17_n_2762 = ~(mul_34_17_n_1704 | mul_34_17_n_402);
 assign mul_34_17_n_2761 = ~(mul_34_17_n_1728 | mul_34_17_n_403);
 assign mul_34_17_n_2760 = ~(mul_34_17_n_1708 | mul_34_17_n_419);
 assign mul_34_17_n_2759 = ~(mul_34_17_n_1731 | mul_34_17_n_404);
 assign mul_34_17_n_2758 = ~(mul_34_17_n_1705 | mul_34_17_n_405);
 assign mul_34_17_n_2757 = ~(mul_34_17_n_1726 | mul_34_17_n_406);
 assign mul_34_17_n_2756 = ~(mul_34_17_n_1722 | mul_34_17_n_420);
 assign mul_34_17_n_2755 = ~(mul_34_17_n_1712 | mul_34_17_n_407);
 assign mul_34_17_n_2754 = ~(mul_34_17_n_1750 | mul_34_17_n_2577);
 assign mul_34_17_n_2711 = ~(mul_34_17_n_1713 | mul_34_17_n_409);
 assign mul_34_17_n_2710 = ~(mul_34_17_n_1699 | mul_34_17_n_422);
 assign mul_34_17_n_2709 = ~(mul_34_17_n_1720 | mul_34_17_n_423);
 assign mul_34_17_n_2708 = ~(mul_34_17_n_1727 | mul_34_17_n_410);
 assign mul_34_17_n_2707 = ~(mul_34_17_n_1714 | mul_34_17_n_424);
 assign mul_34_17_n_2706 = ~(mul_34_17_n_1707 | mul_34_17_n_425);
 assign mul_34_17_n_2705 = ~(mul_34_17_n_1732 | mul_34_17_n_408);
 assign mul_34_17_n_2704 = ~(mul_34_17_n_1709 | mul_34_17_n_421);
 assign mul_34_17_n_2703 = ~(mul_34_17_n_675 & mul_34_17_n_981);
 assign mul_34_17_n_2753 = ~(mul_34_17_n_680 | mul_34_17_n_875);
 assign mul_34_17_n_2752 = ~(mul_34_17_n_666 | mul_34_17_n_1219);
 assign mul_34_17_n_2751 = ~(mul_34_17_n_1736 | mul_34_17_n_2698);
 assign mul_34_17_n_2750 = ~(mul_34_17_n_668 | mul_34_17_n_1154);
 assign mul_34_17_n_2749 = ~(mul_34_17_n_658 | mul_34_17_n_1498);
 assign mul_34_17_n_2748 = ~(mul_34_17_n_668 | mul_34_17_n_1181);
 assign mul_34_17_n_2747 = ~(mul_34_17_n_654 | mul_34_17_n_1657);
 assign mul_34_17_n_2746 = ~(mul_34_17_n_659 & mul_34_17_n_1480);
 assign mul_34_17_n_2745 = ~(mul_34_17_n_689 & mul_34_17_n_756);
 assign mul_34_17_n_2744 = ~(mul_34_17_n_1744 | mul_34_17_n_2289);
 assign mul_34_17_n_2702 = ~(mul_34_17_n_657 & mul_34_17_n_1560);
 assign mul_34_17_n_2743 = ~(mul_34_17_n_1744 | mul_34_17_n_411);
 assign mul_34_17_n_2742 = ~(mul_34_17_n_683 & {in1[0]});
 assign mul_34_17_n_2741 = ~(mul_34_17_n_1735 & {in1[0]});
 assign mul_34_17_n_2740 = ~(mul_34_17_n_1749 & {in1[0]});
 assign mul_34_17_n_2739 = ~(mul_34_17_n_1753 & {in1[0]});
 assign mul_34_17_n_2738 = ~(mul_34_17_n_684 | mul_34_17_n_411);
 assign mul_34_17_n_2737 = ~(mul_34_17_n_667 & {in1[0]});
 assign mul_34_17_n_2736 = ~(mul_34_17_n_1739 & {in1[0]});
 assign mul_34_17_n_2735 = ~(mul_34_17_n_657 & {in1[0]});
 assign mul_34_17_n_2734 = ~(mul_34_17_n_681 & {in1[0]});
 assign mul_34_17_n_2733 = ~(mul_34_17_n_665 & {in1[0]});
 assign mul_34_17_n_2732 = ~(mul_34_17_n_679 & {in1[0]});
 assign mul_34_17_n_2731 = ~(mul_34_17_n_691 & {in1[0]});
 assign mul_34_17_n_2730 = ~(mul_34_17_n_1737 & {in1[0]});
 assign mul_34_17_n_2729 = ~(mul_34_17_n_689 & {in1[0]});
 assign mul_34_17_n_2728 = ~(mul_34_17_n_671 & {in1[0]});
 assign mul_34_17_n_2727 = ~(mul_34_17_n_1757 & {in1[0]});
 assign mul_34_17_n_2726 = ~(mul_34_17_n_669 & {in1[0]});
 assign mul_34_17_n_2725 = ~(mul_34_17_n_655 & {in1[0]});
 assign mul_34_17_n_2724 = ~(mul_34_17_n_677 & {in1[0]});
 assign mul_34_17_n_2723 = ~(mul_34_17_n_1755 & {in1[0]});
 assign mul_34_17_n_2722 = ~(mul_34_17_n_1742 | mul_34_17_n_411);
 assign mul_34_17_n_2721 = ~(mul_34_17_n_675 & {in1[0]});
 assign mul_34_17_n_2720 = ~(mul_34_17_n_1747 & {in1[0]});
 assign mul_34_17_n_2719 = ~(mul_34_17_n_1751 & {in1[0]});
 assign mul_34_17_n_2718 = ~(mul_34_17_n_659 & {in1[0]});
 assign mul_34_17_n_2717 = ~(mul_34_17_n_687 & {in1[0]});
 assign mul_34_17_n_2716 = ~(mul_34_17_n_673 & {in1[0]});
 assign mul_34_17_n_2715 = ~(mul_34_17_n_661 & {in1[0]});
 assign mul_34_17_n_2714 = ~(mul_34_17_n_1741 & {in1[0]});
 assign mul_34_17_n_2713 = ~(mul_34_17_n_663 & {in1[0]});
 assign mul_34_17_n_2712 = ((mul_34_17_n_516 | {in2[0]}) & (mul_34_17_n_485 | mul_34_17_n_486));
 assign mul_34_17_n_2700 = ~mul_34_17_n_2699;
 assign mul_34_17_n_2698 = ~mul_34_17_n_2697;
 assign mul_34_17_n_2679 = ~mul_34_17_n_2678;
 assign mul_34_17_n_2672 = ~mul_34_17_n_2671;
 assign mul_34_17_n_2661 = ~mul_34_17_n_2660;
 assign mul_34_17_n_2657 = ~mul_34_17_n_2656;
 assign mul_34_17_n_2653 = ~mul_34_17_n_2652;
 assign mul_34_17_n_2642 = ~mul_34_17_n_2641;
 assign mul_34_17_n_2637 = ~mul_34_17_n_2636;
 assign mul_34_17_n_2630 = ~mul_34_17_n_2629;
 assign mul_34_17_n_2625 = ~mul_34_17_n_2624;
 assign mul_34_17_n_2620 = ~mul_34_17_n_2619;
 assign mul_34_17_n_2615 = ~mul_34_17_n_2614;
 assign mul_34_17_n_2602 = ~mul_34_17_n_2601;
 assign mul_34_17_n_2599 = ~mul_34_17_n_2598;
 assign mul_34_17_n_2596 = ~mul_34_17_n_2595;
 assign mul_34_17_n_2584 = ~mul_34_17_n_2583;
 assign mul_34_17_n_2582 = ~mul_34_17_n_2581;
 assign mul_34_17_n_2578 = ~mul_34_17_n_2577;
 assign mul_34_17_n_2575 = ~mul_34_17_n_2574;
 assign mul_34_17_n_2572 = ~mul_34_17_n_2571;
 assign mul_34_17_n_2564 = ~mul_34_17_n_2563;
 assign mul_34_17_n_2559 = ~mul_34_17_n_2558;
 assign mul_34_17_n_2554 = ~mul_34_17_n_2553;
 assign mul_34_17_n_2552 = ~mul_34_17_n_2551;
 assign mul_34_17_n_2540 = ~mul_34_17_n_2539;
 assign mul_34_17_n_2534 = ~mul_34_17_n_2533;
 assign mul_34_17_n_2530 = ~mul_34_17_n_2529;
 assign mul_34_17_n_2527 = ~mul_34_17_n_2526;
 assign mul_34_17_n_2523 = ~mul_34_17_n_2522;
 assign mul_34_17_n_2521 = ~mul_34_17_n_2520;
 assign mul_34_17_n_2517 = ~mul_34_17_n_2516;
 assign mul_34_17_n_2515 = ~mul_34_17_n_2514;
 assign mul_34_17_n_2513 = ~mul_34_17_n_2512;
 assign mul_34_17_n_2507 = ~mul_34_17_n_2506;
 assign mul_34_17_n_2493 = ~mul_34_17_n_2492;
 assign mul_34_17_n_2490 = ~mul_34_17_n_2489;
 assign mul_34_17_n_2486 = ~mul_34_17_n_2485;
 assign mul_34_17_n_2481 = ~mul_34_17_n_2480;
 assign mul_34_17_n_2478 = ~mul_34_17_n_2477;
 assign mul_34_17_n_2475 = ~mul_34_17_n_2474;
 assign mul_34_17_n_2470 = ~mul_34_17_n_2469;
 assign mul_34_17_n_2467 = ~mul_34_17_n_2466;
 assign mul_34_17_n_2465 = ~mul_34_17_n_2464;
 assign mul_34_17_n_2457 = ~mul_34_17_n_2456;
 assign mul_34_17_n_2450 = ~mul_34_17_n_2449;
 assign mul_34_17_n_2446 = ~mul_34_17_n_2445;
 assign mul_34_17_n_2443 = ~mul_34_17_n_2442;
 assign mul_34_17_n_2440 = ~mul_34_17_n_2439;
 assign mul_34_17_n_2431 = ~mul_34_17_n_2430;
 assign mul_34_17_n_2425 = ~mul_34_17_n_2424;
 assign mul_34_17_n_2422 = ~mul_34_17_n_2421;
 assign mul_34_17_n_2417 = ~mul_34_17_n_2416;
 assign mul_34_17_n_2409 = ~mul_34_17_n_2408;
 assign mul_34_17_n_2406 = ~mul_34_17_n_2405;
 assign mul_34_17_n_2394 = ~mul_34_17_n_2393;
 assign mul_34_17_n_2388 = ~mul_34_17_n_2387;
 assign mul_34_17_n_2384 = ~mul_34_17_n_2383;
 assign mul_34_17_n_2375 = ~mul_34_17_n_2374;
 assign mul_34_17_n_2373 = ~mul_34_17_n_2372;
 assign mul_34_17_n_2365 = ~mul_34_17_n_2364;
 assign mul_34_17_n_2361 = ~mul_34_17_n_2360;
 assign mul_34_17_n_2358 = ~mul_34_17_n_2357;
 assign mul_34_17_n_2352 = ~mul_34_17_n_2351;
 assign mul_34_17_n_2350 = ~mul_34_17_n_2349;
 assign mul_34_17_n_2343 = ~mul_34_17_n_2342;
 assign mul_34_17_n_2328 = ~mul_34_17_n_2327;
 assign mul_34_17_n_2326 = ~mul_34_17_n_2325;
 assign mul_34_17_n_2324 = ~mul_34_17_n_2323;
 assign mul_34_17_n_2318 = ~mul_34_17_n_2317;
 assign mul_34_17_n_2316 = ~mul_34_17_n_2315;
 assign mul_34_17_n_2314 = ~mul_34_17_n_2313;
 assign mul_34_17_n_2311 = ~mul_34_17_n_2310;
 assign mul_34_17_n_2307 = ~mul_34_17_n_2306;
 assign mul_34_17_n_2305 = ~mul_34_17_n_2304;
 assign mul_34_17_n_2295 = ~mul_34_17_n_2294;
 assign mul_34_17_n_2292 = ~mul_34_17_n_2291;
 assign mul_34_17_n_2290 = ~mul_34_17_n_2289;
 assign mul_34_17_n_2287 = ~mul_34_17_n_2286;
 assign mul_34_17_n_2281 = ~mul_34_17_n_2280;
 assign mul_34_17_n_2278 = ~mul_34_17_n_2277;
 assign mul_34_17_n_2272 = ~mul_34_17_n_2271;
 assign mul_34_17_n_2270 = ~mul_34_17_n_2269;
 assign mul_34_17_n_2266 = ~mul_34_17_n_2265;
 assign mul_34_17_n_2257 = ~mul_34_17_n_2256;
 assign mul_34_17_n_2254 = ~mul_34_17_n_2253;
 assign mul_34_17_n_2251 = ~mul_34_17_n_2250;
 assign mul_34_17_n_2249 = ~mul_34_17_n_2248;
 assign mul_34_17_n_2243 = ~mul_34_17_n_2242;
 assign mul_34_17_n_2233 = ~mul_34_17_n_2232;
 assign mul_34_17_n_2225 = ~mul_34_17_n_2224;
 assign mul_34_17_n_2202 = ~mul_34_17_n_2201;
 assign mul_34_17_n_2198 = ~mul_34_17_n_2197;
 assign mul_34_17_n_2182 = ~mul_34_17_n_2181;
 assign mul_34_17_n_2180 = ~mul_34_17_n_2179;
 assign mul_34_17_n_2177 = ~mul_34_17_n_2176;
 assign mul_34_17_n_2169 = ~mul_34_17_n_2168;
 assign mul_34_17_n_2165 = ~mul_34_17_n_2164;
 assign mul_34_17_n_2162 = ~mul_34_17_n_2161;
 assign mul_34_17_n_2158 = ~mul_34_17_n_2157;
 assign mul_34_17_n_2153 = ~mul_34_17_n_2152;
 assign mul_34_17_n_2143 = ~mul_34_17_n_2142;
 assign mul_34_17_n_2140 = ~mul_34_17_n_2139;
 assign mul_34_17_n_2137 = ~mul_34_17_n_2136;
 assign mul_34_17_n_2128 = ~mul_34_17_n_2127;
 assign mul_34_17_n_2126 = ~mul_34_17_n_2125;
 assign mul_34_17_n_2122 = ~mul_34_17_n_2121;
 assign mul_34_17_n_2117 = ~mul_34_17_n_2116;
 assign mul_34_17_n_2113 = ~mul_34_17_n_2112;
 assign mul_34_17_n_2106 = ~mul_34_17_n_2105;
 assign mul_34_17_n_2104 = ~mul_34_17_n_2103;
 assign mul_34_17_n_2097 = ~mul_34_17_n_2096;
 assign mul_34_17_n_2094 = ~mul_34_17_n_2093;
 assign mul_34_17_n_2092 = ~mul_34_17_n_2091;
 assign mul_34_17_n_2086 = ~mul_34_17_n_2085;
 assign mul_34_17_n_2081 = ~mul_34_17_n_2080;
 assign mul_34_17_n_2078 = ~mul_34_17_n_2077;
 assign mul_34_17_n_2075 = ~mul_34_17_n_2074;
 assign mul_34_17_n_2073 = ~mul_34_17_n_2072;
 assign mul_34_17_n_2069 = ~mul_34_17_n_2068;
 assign mul_34_17_n_2065 = ~mul_34_17_n_2064;
 assign mul_34_17_n_2062 = ~mul_34_17_n_2061;
 assign mul_34_17_n_2051 = ~mul_34_17_n_2050;
 assign mul_34_17_n_2046 = ~mul_34_17_n_2045;
 assign mul_34_17_n_2041 = ~mul_34_17_n_2040;
 assign mul_34_17_n_2035 = ~mul_34_17_n_2034;
 assign mul_34_17_n_2033 = ~mul_34_17_n_2032;
 assign mul_34_17_n_2027 = ~mul_34_17_n_2026;
 assign mul_34_17_n_2025 = ~mul_34_17_n_2024;
 assign mul_34_17_n_2023 = ~mul_34_17_n_2022;
 assign mul_34_17_n_2021 = ~mul_34_17_n_2020;
 assign mul_34_17_n_2017 = ~mul_34_17_n_2016;
 assign mul_34_17_n_2014 = ~mul_34_17_n_2013;
 assign mul_34_17_n_2010 = ~mul_34_17_n_2009;
 assign mul_34_17_n_2002 = ~mul_34_17_n_2001;
 assign mul_34_17_n_2000 = ~mul_34_17_n_1999;
 assign mul_34_17_n_1987 = ~mul_34_17_n_1986;
 assign mul_34_17_n_1985 = ~mul_34_17_n_1984;
 assign mul_34_17_n_1982 = ~mul_34_17_n_1981;
 assign mul_34_17_n_1980 = ~mul_34_17_n_1979;
 assign mul_34_17_n_1977 = ~mul_34_17_n_1976;
 assign mul_34_17_n_1975 = ~mul_34_17_n_1974;
 assign mul_34_17_n_1970 = ~mul_34_17_n_1969;
 assign mul_34_17_n_1966 = ~mul_34_17_n_1965;
 assign mul_34_17_n_1964 = ~mul_34_17_n_1963;
 assign mul_34_17_n_1959 = ~mul_34_17_n_1958;
 assign mul_34_17_n_1953 = ~mul_34_17_n_1952;
 assign mul_34_17_n_1951 = ~mul_34_17_n_1950;
 assign mul_34_17_n_1949 = ~mul_34_17_n_1948;
 assign mul_34_17_n_1942 = ~mul_34_17_n_1941;
 assign mul_34_17_n_1939 = ~mul_34_17_n_1938;
 assign mul_34_17_n_1936 = ~mul_34_17_n_1935;
 assign mul_34_17_n_1924 = ~mul_34_17_n_1923;
 assign mul_34_17_n_1920 = ~mul_34_17_n_1919;
 assign mul_34_17_n_1915 = ~mul_34_17_n_1914;
 assign mul_34_17_n_1905 = ~mul_34_17_n_1904;
 assign mul_34_17_n_1901 = ~mul_34_17_n_1900;
 assign mul_34_17_n_1899 = ~mul_34_17_n_1898;
 assign mul_34_17_n_1897 = ~mul_34_17_n_1896;
 assign mul_34_17_n_1888 = ~mul_34_17_n_1887;
 assign mul_34_17_n_1885 = ~mul_34_17_n_1884;
 assign mul_34_17_n_1882 = ~mul_34_17_n_1881;
 assign mul_34_17_n_1880 = ~mul_34_17_n_1879;
 assign mul_34_17_n_1868 = ~mul_34_17_n_1867;
 assign mul_34_17_n_1865 = ~mul_34_17_n_1864;
 assign mul_34_17_n_1862 = ~mul_34_17_n_1861;
 assign mul_34_17_n_1845 = ~mul_34_17_n_1844;
 assign mul_34_17_n_1843 = ~mul_34_17_n_1842;
 assign mul_34_17_n_1773 = ~mul_34_17_n_1772;
 assign mul_34_17_n_1769 = ~mul_34_17_n_1768;
 assign mul_34_17_n_1767 = ~mul_34_17_n_1766;
 assign mul_34_17_n_1762 = ~mul_34_17_n_1761;
 assign mul_34_17_n_1756 = ~mul_34_17_n_1757;
 assign mul_34_17_n_1754 = ~mul_34_17_n_1755;
 assign mul_34_17_n_1752 = ~mul_34_17_n_1753;
 assign mul_34_17_n_1750 = ~mul_34_17_n_1751;
 assign mul_34_17_n_1748 = ~mul_34_17_n_1749;
 assign mul_34_17_n_1746 = ~mul_34_17_n_1747;
 assign mul_34_17_n_1744 = ~mul_34_17_n_1745;
 assign mul_34_17_n_1742 = ~mul_34_17_n_1743;
 assign mul_34_17_n_1740 = ~mul_34_17_n_1741;
 assign mul_34_17_n_1738 = ~mul_34_17_n_1739;
 assign mul_34_17_n_1736 = ~mul_34_17_n_1737;
 assign mul_34_17_n_1734 = ~mul_34_17_n_1735;
 assign mul_34_17_n_1733 = ~(mul_34_17_n_542 | mul_34_17_n_414);
 assign mul_34_17_n_1732 = ~(mul_34_17_n_568 | mul_34_17_n_421);
 assign mul_34_17_n_1731 = ~(mul_34_17_n_548 | mul_34_17_n_419);
 assign mul_34_17_n_1730 = ~(mul_34_17_n_555 | mul_34_17_n_416);
 assign mul_34_17_n_1729 = ~(mul_34_17_n_559 | mul_34_17_n_418);
 assign mul_34_17_n_1728 = ~(mul_34_17_n_552 | mul_34_17_n_402);
 assign mul_34_17_n_1727 = ~(mul_34_17_n_540 | mul_34_17_n_423);
 assign mul_34_17_n_1726 = ~(mul_34_17_n_562 | mul_34_17_n_405);
 assign mul_34_17_n_1725 = ~(mul_34_17_n_549 | mul_34_17_n_417);
 assign mul_34_17_n_1724 = ~(mul_34_17_n_547 | mul_34_17_n_395);
 assign mul_34_17_n_1723 = ~(mul_34_17_n_560 | mul_34_17_n_398);
 assign mul_34_17_n_1722 = ~(mul_34_17_n_496 | mul_34_17_n_406);
 assign mul_34_17_n_1721 = ~(mul_34_17_n_567 | mul_34_17_n_399);
 assign mul_34_17_n_1720 = ~(mul_34_17_n_571 | mul_34_17_n_422);
 assign mul_34_17_n_1719 = ~(mul_34_17_n_508 | mul_34_17_n_394);
 assign mul_34_17_n_1718 = ~(mul_34_17_n_531 | mul_34_17_n_397);
 assign mul_34_17_n_1717 = ~(mul_34_17_n_495 | mul_34_17_n_412);
 assign mul_34_17_n_1716 = ~(mul_34_17_n_532 | mul_34_17_n_393);
 assign mul_34_17_n_1715 = ~(mul_34_17_n_476 | mul_34_17_n_413);
 assign mul_34_17_n_1714 = ~(mul_34_17_n_509 | mul_34_17_n_410);
 assign mul_34_17_n_1713 = ~(mul_34_17_n_538 | mul_34_17_n_408);
 assign mul_34_17_n_1712 = ~(mul_34_17_n_513 | mul_34_17_n_420);
 assign mul_34_17_n_1711 = ~(mul_34_17_n_536 | mul_34_17_n_396);
 assign mul_34_17_n_1710 = ~(mul_34_17_n_544 | mul_34_17_n_400);
 assign mul_34_17_n_1709 = ~(mul_34_17_n_566 | mul_34_17_n_407);
 assign mul_34_17_n_1708 = ~(mul_34_17_n_512 | mul_34_17_n_403);
 assign mul_34_17_n_1707 = ~(mul_34_17_n_504 | mul_34_17_n_424);
 assign mul_34_17_n_1706 = ~(mul_34_17_n_511 | mul_34_17_n_415);
 assign mul_34_17_n_1705 = ~(mul_34_17_n_497 | mul_34_17_n_404);
 assign mul_34_17_n_1704 = ~(mul_34_17_n_564 | mul_34_17_n_401);
 assign mul_34_17_n_1703 = ({in2[1]} ^ {in1[0]});
 assign mul_34_17_n_1702 = ~({in2[61]} ^ {in1[0]});
 assign mul_34_17_n_1701 = ~({in2[55]} ^ {in1[0]});
 assign mul_34_17_n_1700 = ({in2[23]} ^ {in1[63]});
 assign mul_34_17_n_1699 = ~(mul_34_17_n_551 | mul_34_17_n_409);
 assign mul_34_17_n_2701 = ~({in2[19]} ^ {in1[23]});
 assign mul_34_17_n_2699 = ~({in2[17]} ^ {in1[9]});
 assign mul_34_17_n_2697 = ({in2[13]} ^ {in1[42]});
 assign mul_34_17_n_2696 = ~({in2[5]} ^ {in1[23]});
 assign mul_34_17_n_2695 = ({in2[15]} ^ {in1[43]});
 assign mul_34_17_n_2694 = ({in2[19]} ^ {in1[62]});
 assign mul_34_17_n_2693 = ~({in2[3]} ^ {in1[59]});
 assign mul_34_17_n_2692 = ~({in2[19]} ^ {in1[11]});
 assign mul_34_17_n_2691 = ({in2[5]} ^ {in1[47]});
 assign mul_34_17_n_2690 = ({in2[19]} ^ {in1[35]});
 assign mul_34_17_n_2689 = ({in2[3]} ^ {in1[2]});
 assign mul_34_17_n_2688 = ~({in2[19]} ^ {in1[43]});
 assign mul_34_17_n_2687 = ({in2[11]} ^ {in1[24]});
 assign mul_34_17_n_2686 = ({in2[3]} ^ {in1[5]});
 assign mul_34_17_n_2685 = ~({in2[11]} ^ {in1[14]});
 assign mul_34_17_n_2684 = ({in2[7]} ^ {in1[5]});
 assign mul_34_17_n_2683 = ~({in2[19]} ^ {in1[42]});
 assign mul_34_17_n_2682 = ({in2[3]} ^ {in1[52]});
 assign mul_34_17_n_2681 = ~({in2[23]} ^ {in1[42]});
 assign mul_34_17_n_2680 = ({in2[21]} ^ {in1[35]});
 assign mul_34_17_n_2678 = ~({in2[9]} ^ {in1[22]});
 assign mul_34_17_n_2677 = ~({in2[21]} ^ {in1[6]});
 assign mul_34_17_n_2676 = ({in2[23]} ^ {in1[12]});
 assign mul_34_17_n_2675 = ~({in2[9]} ^ {in1[59]});
 assign mul_34_17_n_2674 = ~({in2[13]} ^ {in1[36]});
 assign mul_34_17_n_2673 = ({in2[17]} ^ {in1[47]});
 assign mul_34_17_n_2671 = ~({in2[7]} ^ {in1[33]});
 assign mul_34_17_n_2670 = ({in2[23]} ^ {in1[61]});
 assign mul_34_17_n_2669 = ({in2[9]} ^ {in1[11]});
 assign mul_34_17_n_2668 = ({in2[23]} ^ {in1[6]});
 assign mul_34_17_n_2667 = ({in2[23]} ^ {in1[35]});
 assign mul_34_17_n_2666 = ({in2[11]} ^ {in1[45]});
 assign mul_34_17_n_2665 = ({in2[7]} ^ {in1[42]});
 assign mul_34_17_n_2664 = ({in2[15]} ^ {in1[39]});
 assign mul_34_17_n_2663 = ~({in2[5]} ^ {in1[12]});
 assign mul_34_17_n_2662 = ({in2[23]} ^ {in1[7]});
 assign mul_34_17_n_2660 = ~({in2[17]} ^ {in1[3]});
 assign mul_34_17_n_2659 = ({in2[19]} ^ {in1[38]});
 assign mul_34_17_n_2658 = ({in2[25]} ^ {in1[1]});
 assign mul_34_17_n_2656 = ~({in2[23]} ^ {in1[1]});
 assign mul_34_17_n_2655 = ({in2[11]} ^ {in1[44]});
 assign mul_34_17_n_2654 = ({in2[9]} ^ {in1[12]});
 assign mul_34_17_n_2652 = ~({in2[13]} ^ {in1[16]});
 assign mul_34_17_n_2651 = ({in2[3]} ^ {in1[31]});
 assign mul_34_17_n_2650 = ~({in2[21]} ^ {in1[25]});
 assign mul_34_17_n_2649 = ({in2[23]} ^ {in1[62]});
 assign mul_34_17_n_2648 = ({in2[15]} ^ {in1[50]});
 assign mul_34_17_n_2647 = ({in2[5]} ^ {in1[59]});
 assign mul_34_17_n_2646 = ~({in2[19]} ^ {in1[13]});
 assign mul_34_17_n_2645 = ~({in2[7]} ^ {in1[62]});
 assign mul_34_17_n_2644 = ({in2[9]} ^ {in1[48]});
 assign mul_34_17_n_2643 = ({in2[3]} ^ {in1[46]});
 assign mul_34_17_n_2641 = ~({in2[3]} ^ {in1[12]});
 assign mul_34_17_n_2640 = ~({in2[9]} ^ {in1[35]});
 assign mul_34_17_n_2639 = ({in2[11]} ^ {in1[50]});
 assign mul_34_17_n_2638 = ({in2[5]} ^ {in1[45]});
 assign mul_34_17_n_1698 = ~(mul_34_17_n_523 | mul_34_17_n_526);
 assign mul_34_17_n_2636 = ({in2[3]} ^ {in1[17]});
 assign mul_34_17_n_2635 = ({in2[9]} ^ {in1[21]});
 assign mul_34_17_n_2634 = ~({in2[15]} ^ {in1[34]});
 assign mul_34_17_n_2633 = ~({in2[19]} ^ {in1[55]});
 assign mul_34_17_n_2632 = ({in2[17]} ^ {in1[40]});
 assign mul_34_17_n_2631 = ({in2[13]} ^ {in1[44]});
 assign mul_34_17_n_2629 = ~({in2[19]} ^ {in1[61]});
 assign mul_34_17_n_2628 = ~({in2[23]} ^ {in1[27]});
 assign mul_34_17_n_2627 = ({in2[13]} ^ {in1[14]});
 assign mul_34_17_n_2626 = ({in2[9]} ^ {in1[26]});
 assign mul_34_17_n_2624 = ~({in2[11]} ^ {in1[59]});
 assign mul_34_17_n_2623 = ({in2[9]} ^ {in1[45]});
 assign mul_34_17_n_2622 = ({in2[21]} ^ {in1[30]});
 assign mul_34_17_n_2621 = ({in2[17]} ^ {in1[19]});
 assign mul_34_17_n_2619 = ~({in2[21]} ^ {in1[47]});
 assign mul_34_17_n_2618 = ({in2[13]} ^ {in1[1]});
 assign mul_34_17_n_2617 = ({in2[5]} ^ {in1[25]});
 assign mul_34_17_n_2616 = ({in2[17]} ^ {in1[4]});
 assign mul_34_17_n_2614 = ~({in2[25]} ^ {in1[35]});
 assign mul_34_17_n_2613 = ~({in2[15]} ^ {in1[9]});
 assign mul_34_17_n_2612 = ({in2[15]} ^ {in1[46]});
 assign mul_34_17_n_2611 = ({in2[13]} ^ {in1[54]});
 assign mul_34_17_n_2610 = ~({in2[23]} ^ {in1[26]});
 assign mul_34_17_n_2609 = ({in2[15]} ^ {in1[47]});
 assign mul_34_17_n_2608 = ~({in2[23]} ^ {in1[24]});
 assign mul_34_17_n_2607 = ~({in2[19]} ^ {in1[30]});
 assign mul_34_17_n_2606 = ~({in2[9]} ^ {in1[2]});
 assign mul_34_17_n_2605 = ~({in2[21]} ^ {in1[3]});
 assign mul_34_17_n_2604 = ({in2[7]} ^ {in1[51]});
 assign mul_34_17_n_2603 = ~({in2[9]} ^ {in1[36]});
 assign mul_34_17_n_2601 = ~({in2[19]} ^ {in1[60]});
 assign mul_34_17_n_2600 = ~({in2[17]} ^ {in1[62]});
 assign mul_34_17_n_2598 = ~({in2[9]} ^ {in1[10]});
 assign mul_34_17_n_1697 = ({in2[21]} ^ {in1[63]});
 assign mul_34_17_n_2597 = ({in2[3]} ^ {in1[57]});
 assign mul_34_17_n_2595 = ~({in2[11]} ^ {in1[54]});
 assign mul_34_17_n_2594 = ({in2[21]} ^ {in1[13]});
 assign mul_34_17_n_2593 = ({in2[21]} ^ {in1[58]});
 assign mul_34_17_n_2592 = ~({in2[15]} ^ {in1[56]});
 assign mul_34_17_n_2591 = ({in2[19]} ^ {in1[15]});
 assign mul_34_17_n_2590 = ({in2[21]} ^ {in1[44]});
 assign mul_34_17_n_2589 = ({in2[17]} ^ {in1[12]});
 assign mul_34_17_n_2588 = ({in2[23]} ^ {in1[13]});
 assign mul_34_17_n_2587 = ({in2[3]} ^ {in1[50]});
 assign mul_34_17_n_2586 = ({in2[11]} ^ {in1[40]});
 assign mul_34_17_n_2585 = ~({in2[5]} ^ {in1[13]});
 assign mul_34_17_n_2583 = ~({in2[9]} ^ {in1[23]});
 assign mul_34_17_n_2581 = ({in2[9]} ^ {in1[13]});
 assign mul_34_17_n_2580 = ({in2[9]} ^ {in1[27]});
 assign mul_34_17_n_2579 = ({in2[11]} ^ {in1[17]});
 assign mul_34_17_n_2577 = ~({in2[9]} ^ {in1[44]});
 assign mul_34_17_n_2576 = ({in2[7]} ^ {in1[60]});
 assign mul_34_17_n_2574 = ~({in2[7]} ^ {in1[61]});
 assign mul_34_17_n_2573 = ({in2[13]} ^ {in1[18]});
 assign mul_34_17_n_2571 = ~({in2[11]} ^ {in1[34]});
 assign mul_34_17_n_2570 = ({in2[5]} ^ {in1[29]});
 assign mul_34_17_n_2569 = ({in2[7]} ^ {in1[47]});
 assign mul_34_17_n_2568 = ({in2[17]} ^ {in1[43]});
 assign mul_34_17_n_2567 = ({in2[21]} ^ {in1[11]});
 assign mul_34_17_n_2566 = ~({in2[15]} ^ {in1[8]});
 assign mul_34_17_n_2565 = ({in2[19]} ^ {in1[17]});
 assign mul_34_17_n_2563 = ~({in2[11]} ^ {in1[48]});
 assign mul_34_17_n_2562 = ({in2[5]} ^ {in1[9]});
 assign mul_34_17_n_2561 = ({in2[3]} ^ {in1[26]});
 assign mul_34_17_n_2560 = ~({in2[5]} ^ {in1[4]});
 assign mul_34_17_n_2558 = ({in2[9]} ^ {in1[28]});
 assign mul_34_17_n_2557 = ({in2[23]} ^ {in1[55]});
 assign mul_34_17_n_2556 = ~({in2[7]} ^ {in1[20]});
 assign mul_34_17_n_2555 = ~({in2[9]} ^ {in1[18]});
 assign mul_34_17_n_2553 = ({in2[13]} ^ {in1[10]});
 assign mul_34_17_n_2551 = ~({in2[13]} ^ {in1[45]});
 assign mul_34_17_n_2550 = ~({in2[13]} ^ {in1[11]});
 assign mul_34_17_n_2549 = ~({in2[7]} ^ {in1[22]});
 assign mul_34_17_n_2548 = ~({in2[23]} ^ {in1[41]});
 assign mul_34_17_n_2547 = ({in2[23]} ^ {in1[11]});
 assign mul_34_17_n_2546 = ({in2[13]} ^ {in1[40]});
 assign mul_34_17_n_2545 = ({in2[3]} ^ {in1[11]});
 assign mul_34_17_n_2544 = ({in2[13]} ^ {in1[49]});
 assign mul_34_17_n_2543 = ({in2[11]} ^ {in1[56]});
 assign mul_34_17_n_2542 = ({in2[25]} ^ {in1[48]});
 assign mul_34_17_n_2541 = ({in2[17]} ^ {in1[13]});
 assign mul_34_17_n_2539 = ~({in2[21]} ^ {in1[20]});
 assign mul_34_17_n_2538 = ~({in2[7]} ^ {in1[17]});
 assign mul_34_17_n_2537 = ~({in2[17]} ^ {in1[2]});
 assign mul_34_17_n_2536 = ~({in2[13]} ^ {in1[28]});
 assign mul_34_17_n_2535 = ({in2[15]} ^ {in1[42]});
 assign mul_34_17_n_1696 = ~(mul_34_17_n_527 | mul_34_17_n_528);
 assign mul_34_17_n_2533 = ~({in2[7]} ^ {in1[58]});
 assign mul_34_17_n_2532 = ({in2[7]} ^ {in1[28]});
 assign mul_34_17_n_2531 = ~({in2[9]} ^ {in1[15]});
 assign mul_34_17_n_2529 = ~({in2[3]} ^ {in1[37]});
 assign mul_34_17_n_2528 = ({in2[19]} ^ {in1[33]});
 assign mul_34_17_n_2526 = ~({in2[9]} ^ {in1[32]});
 assign mul_34_17_n_2525 = ~({in2[13]} ^ {in1[30]});
 assign mul_34_17_n_2524 = ({in2[21]} ^ {in1[1]});
 assign mul_34_17_n_2522 = ({in2[13]} ^ {in1[39]});
 assign mul_34_17_n_2520 = ~({in2[19]} ^ {in1[18]});
 assign mul_34_17_n_2519 = ~({in2[5]} ^ {in1[39]});
 assign mul_34_17_n_2518 = ({in2[3]} ^ {in1[28]});
 assign mul_34_17_n_2516 = ~({in2[19]} ^ {in1[45]});
 assign mul_34_17_n_2514 = ~({in2[17]} ^ {in1[49]});
 assign mul_34_17_n_2512 = ~({in2[19]} ^ {in1[47]});
 assign mul_34_17_n_2511 = ~({in2[13]} ^ {in1[59]});
 assign mul_34_17_n_2510 = ~({in2[19]} ^ {in1[6]});
 assign mul_34_17_n_2509 = ~({in2[7]} ^ {in1[54]});
 assign mul_34_17_n_2508 = ~({in2[9]} ^ {in1[37]});
 assign mul_34_17_n_2506 = ~({in2[7]} ^ {in1[40]});
 assign mul_34_17_n_2505 = ({in2[15]} ^ {in1[11]});
 assign mul_34_17_n_2504 = ~({in2[11]} ^ {in1[62]});
 assign mul_34_17_n_2503 = ({in2[13]} ^ {in1[8]});
 assign mul_34_17_n_2502 = ({in2[3]} ^ {in1[53]});
 assign mul_34_17_n_2501 = ({in2[19]} ^ {in1[16]});
 assign mul_34_17_n_2500 = ~({in2[9]} ^ {in1[54]});
 assign mul_34_17_n_2499 = ~({in2[11]} ^ {in1[61]});
 assign mul_34_17_n_2498 = ({in2[21]} ^ {in1[39]});
 assign mul_34_17_n_2497 = ({in2[15]} ^ {in1[62]});
 assign mul_34_17_n_2496 = ~({in2[15]} ^ {in1[6]});
 assign mul_34_17_n_2495 = ~({in2[23]} ^ {in1[46]});
 assign mul_34_17_n_2494 = ~({in2[19]} ^ {in1[54]});
 assign mul_34_17_n_2492 = ~({in2[7]} ^ {in1[2]});
 assign mul_34_17_n_2491 = ({in2[11]} ^ {in1[28]});
 assign mul_34_17_n_2489 = ~({in2[15]} ^ {in1[25]});
 assign mul_34_17_n_2488 = ({in2[15]} ^ {in1[41]});
 assign mul_34_17_n_2487 = ~({in2[11]} ^ {in1[58]});
 assign mul_34_17_n_2485 = ~({in2[7]} ^ {in1[39]});
 assign mul_34_17_n_2484 = ({in2[17]} ^ {in1[44]});
 assign mul_34_17_n_2483 = ({in2[23]} ^ {in1[31]});
 assign mul_34_17_n_2482 = ({in2[3]} ^ {in1[3]});
 assign mul_34_17_n_2480 = ~({in2[3]} ^ {in1[43]});
 assign mul_34_17_n_2479 = ~({in2[15]} ^ {in1[33]});
 assign mul_34_17_n_2477 = ({in2[23]} ^ {in1[15]});
 assign mul_34_17_n_2476 = ({in2[17]} ^ {in1[42]});
 assign mul_34_17_n_2474 = ~({in2[3]} ^ {in1[44]});
 assign mul_34_17_n_2473 = ({in2[17]} ^ {in1[50]});
 assign mul_34_17_n_2472 = ({in2[5]} ^ {in1[61]});
 assign mul_34_17_n_2471 = ~({in2[15]} ^ {in1[31]});
 assign mul_34_17_n_2469 = ~({in2[21]} ^ {in1[41]});
 assign mul_34_17_n_2468 = ({in2[15]} ^ {in1[20]});
 assign mul_34_17_n_2466 = ~({in2[5]} ^ {in1[11]});
 assign mul_34_17_n_2464 = ({in2[13]} ^ {in1[13]});
 assign mul_34_17_n_2463 = ({in2[3]} ^ {in1[62]});
 assign mul_34_17_n_2462 = ~({in2[15]} ^ {in1[7]});
 assign mul_34_17_n_2461 = ({in2[17]} ^ {in1[31]});
 assign mul_34_17_n_2460 = ~({in2[13]} ^ {in1[4]});
 assign mul_34_17_n_2459 = ({in2[9]} ^ {in1[42]});
 assign mul_34_17_n_2458 = ~({in2[11]} ^ {in1[7]});
 assign mul_34_17_n_2456 = ~({in2[9]} ^ {in1[57]});
 assign mul_34_17_n_2455 = ({in2[19]} ^ {in1[32]});
 assign mul_34_17_n_2454 = ({in2[15]} ^ {in1[36]});
 assign mul_34_17_n_2453 = ({in2[5]} ^ {in1[62]});
 assign mul_34_17_n_2452 = ({in2[23]} ^ {in1[44]});
 assign mul_34_17_n_2451 = ({in2[17]} ^ {in1[34]});
 assign mul_34_17_n_2449 = ({in2[15]} ^ {in1[52]});
 assign mul_34_17_n_2448 = ~({in2[9]} ^ {in1[38]});
 assign mul_34_17_n_2447 = ({in2[23]} ^ {in1[29]});
 assign mul_34_17_n_2445 = ~({in2[23]} ^ {in1[23]});
 assign mul_34_17_n_2444 = ({in2[21]} ^ {in1[9]});
 assign mul_34_17_n_2442 = ({in2[17]} ^ {in1[1]});
 assign mul_34_17_n_2441 = ~({in2[19]} ^ {in1[21]});
 assign mul_34_17_n_2439 = ~({in2[5]} ^ {in1[58]});
 assign mul_34_17_n_2438 = ~({in2[17]} ^ {in1[59]});
 assign mul_34_17_n_2437 = ~({in2[9]} ^ {in1[7]});
 assign mul_34_17_n_2436 = ~({in2[13]} ^ {in1[5]});
 assign mul_34_17_n_2435 = ({in2[25]} ^ {in1[11]});
 assign mul_34_17_n_2434 = ({in2[23]} ^ {in1[30]});
 assign mul_34_17_n_2433 = ({in2[21]} ^ {in1[57]});
 assign mul_34_17_n_2432 = ({in2[7]} ^ {in1[50]});
 assign mul_34_17_n_2430 = ~({in2[23]} ^ {in1[53]});
 assign mul_34_17_n_2429 = ({in2[13]} ^ {in1[21]});
 assign mul_34_17_n_2428 = ({in2[21]} ^ {in1[14]});
 assign mul_34_17_n_2427 = ({in2[13]} ^ {in1[23]});
 assign mul_34_17_n_2426 = ({in2[5]} ^ {in1[53]});
 assign mul_34_17_n_2424 = ({in2[15]} ^ {in1[14]});
 assign mul_34_17_n_2423 = ({in2[5]} ^ {in1[34]});
 assign mul_34_17_n_2421 = ~({in2[3]} ^ {in1[42]});
 assign mul_34_17_n_2420 = ~({in2[23]} ^ {in1[50]});
 assign mul_34_17_n_2419 = ~({in2[13]} ^ {in1[31]});
 assign mul_34_17_n_2418 = ({in2[17]} ^ {in1[36]});
 assign mul_34_17_n_2416 = ~({in2[19]} ^ {in1[26]});
 assign mul_34_17_n_2415 = ({in2[7]} ^ {in1[27]});
 assign mul_34_17_n_2414 = ~({in2[19]} ^ {in1[12]});
 assign mul_34_17_n_2413 = ~({in2[9]} ^ {in1[61]});
 assign mul_34_17_n_2412 = ~({in2[5]} ^ {in1[41]});
 assign mul_34_17_n_2411 = ({in2[13]} ^ {in1[26]});
 assign mul_34_17_n_2410 = ~({in2[21]} ^ {in1[26]});
 assign mul_34_17_n_2408 = ~({in2[15]} ^ {in1[12]});
 assign mul_34_17_n_2407 = ~({in2[13]} ^ {in1[38]});
 assign mul_34_17_n_2405 = ~({in2[17]} ^ {in1[48]});
 assign mul_34_17_n_2404 = ({in2[5]} ^ {in1[2]});
 assign mul_34_17_n_2403 = ~({in2[3]} ^ {in1[7]});
 assign mul_34_17_n_2402 = ~({in2[21]} ^ {in1[49]});
 assign mul_34_17_n_2401 = ~({in2[21]} ^ {in1[48]});
 assign mul_34_17_n_2400 = ~({in2[21]} ^ {in1[24]});
 assign mul_34_17_n_2399 = ~({in2[3]} ^ {in1[41]});
 assign mul_34_17_n_2398 = ~({in2[5]} ^ {in1[21]});
 assign mul_34_17_n_2397 = ({in2[21]} ^ {in1[32]});
 assign mul_34_17_n_2396 = ({in2[23]} ^ {in1[10]});
 assign mul_34_17_n_2395 = ({in2[11]} ^ {in1[23]});
 assign mul_34_17_n_2393 = ({in2[13]} ^ {in1[48]});
 assign mul_34_17_n_2392 = ({in2[3]} ^ {in1[24]});
 assign mul_34_17_n_2391 = ({in2[3]} ^ {in1[48]});
 assign mul_34_17_n_1695 = ~(mul_34_17_n_522 | mul_34_17_n_524);
 assign mul_34_17_n_2390 = ({in2[11]} ^ {in1[19]});
 assign mul_34_17_n_2389 = ({in2[11]} ^ {in1[20]});
 assign mul_34_17_n_2387 = ~({in2[9]} ^ {in1[1]});
 assign mul_34_17_n_2386 = ~({in2[17]} ^ {in1[53]});
 assign mul_34_17_n_2385 = ({in2[23]} ^ {in1[52]});
 assign mul_34_17_n_2383 = ~({in2[15]} ^ {in1[35]});
 assign mul_34_17_n_2382 = ({in2[3]} ^ {in1[54]});
 assign mul_34_17_n_2381 = ({in2[5]} ^ {in1[48]});
 assign mul_34_17_n_2380 = ~({in2[13]} ^ {in1[46]});
 assign mul_34_17_n_2379 = ({in2[19]} ^ {in1[34]});
 assign mul_34_17_n_2378 = ({in2[17]} ^ {in1[35]});
 assign mul_34_17_n_2377 = ~({in2[25]} ^ {in1[45]});
 assign mul_34_17_n_2376 = ~({in2[13]} ^ {in1[57]});
 assign mul_34_17_n_2374 = ~({in2[7]} ^ {in1[12]});
 assign mul_34_17_n_2372 = ~({in2[11]} ^ {in1[30]});
 assign mul_34_17_n_2371 = ~({in2[15]} ^ {in1[55]});
 assign mul_34_17_n_2370 = ({in2[15]} ^ {in1[38]});
 assign mul_34_17_n_2369 = ({in2[7]} ^ {in1[57]});
 assign mul_34_17_n_2368 = ~({in2[19]} ^ {in1[24]});
 assign mul_34_17_n_2367 = ~({in2[5]} ^ {in1[14]});
 assign mul_34_17_n_2366 = ({in2[5]} ^ {in1[46]});
 assign mul_34_17_n_2364 = ~({in2[9]} ^ {in1[58]});
 assign mul_34_17_n_2363 = ({in2[17]} ^ {in1[41]});
 assign mul_34_17_n_2362 = ~({in2[9]} ^ {in1[9]});
 assign mul_34_17_n_2360 = ~({in2[3]} ^ {in1[23]});
 assign mul_34_17_n_2359 = ({in2[21]} ^ {in1[43]});
 assign mul_34_17_n_2357 = ~({in2[7]} ^ {in1[8]});
 assign mul_34_17_n_2356 = ~({in2[5]} ^ {in1[55]});
 assign mul_34_17_n_2355 = ({in2[13]} ^ {in1[22]});
 assign mul_34_17_n_2354 = ({in2[11]} ^ {in1[3]});
 assign mul_34_17_n_2353 = ~({in2[21]} ^ {in1[61]});
 assign mul_34_17_n_2351 = ~({in2[11]} ^ {in1[60]});
 assign mul_34_17_n_2349 = ~({in2[9]} ^ {in1[6]});
 assign mul_34_17_n_2348 = ~({in2[15]} ^ {in1[28]});
 assign mul_34_17_n_2347 = ~({in2[13]} ^ {in1[47]});
 assign mul_34_17_n_2346 = ~({in2[13]} ^ {in1[52]});
 assign mul_34_17_n_2345 = ({in2[15]} ^ {in1[37]});
 assign mul_34_17_n_2344 = ({in2[11]} ^ {in1[1]});
 assign mul_34_17_n_2342 = ~({in2[9]} ^ {in1[50]});
 assign mul_34_17_n_2341 = ({in2[7]} ^ {in1[6]});
 assign mul_34_17_n_2340 = ({in2[3]} ^ {in1[25]});
 assign mul_34_17_n_2339 = ({in2[11]} ^ {in1[35]});
 assign mul_34_17_n_2338 = ({in2[21]} ^ {in1[16]});
 assign mul_34_17_n_2337 = ({in2[7]} ^ {in1[31]});
 assign mul_34_17_n_2336 = ~({in2[17]} ^ {in1[27]});
 assign mul_34_17_n_2335 = ~({in2[5]} ^ {in1[22]});
 assign mul_34_17_n_2334 = ({in2[15]} ^ {in1[48]});
 assign mul_34_17_n_2333 = ({in2[15]} ^ {in1[23]});
 assign mul_34_17_n_2332 = ~({in2[13]} ^ {in1[3]});
 assign mul_34_17_n_2331 = ({in2[17]} ^ {in1[17]});
 assign mul_34_17_n_2330 = ~({in2[9]} ^ {in1[19]});
 assign mul_34_17_n_2329 = ~({in2[3]} ^ {in1[15]});
 assign mul_34_17_n_2327 = ~({in2[11]} ^ {in1[4]});
 assign mul_34_17_n_2325 = ~({in2[9]} ^ {in1[43]});
 assign mul_34_17_n_2323 = ({in2[19]} ^ {in1[14]});
 assign mul_34_17_n_2322 = ~({in2[17]} ^ {in1[55]});
 assign mul_34_17_n_2321 = ({in2[15]} ^ {in1[22]});
 assign mul_34_17_n_2320 = ~({in2[5]} ^ {in1[16]});
 assign mul_34_17_n_2319 = ({in2[21]} ^ {in1[38]});
 assign mul_34_17_n_2317 = ~({in2[3]} ^ {in1[33]});
 assign mul_34_17_n_2315 = ~({in2[19]} ^ {in1[40]});
 assign mul_34_17_n_2313 = ~({in2[5]} ^ {in1[35]});
 assign mul_34_17_n_2312 = ({in2[9]} ^ {in1[5]});
 assign mul_34_17_n_2310 = ~({in2[11]} ^ {in1[55]});
 assign mul_34_17_n_2309 = ({in2[11]} ^ {in1[46]});
 assign mul_34_17_n_2308 = ({in2[19]} ^ {in1[48]});
 assign mul_34_17_n_2306 = ({in2[21]} ^ {in1[17]});
 assign mul_34_17_n_2304 = ~({in2[15]} ^ {in1[44]});
 assign mul_34_17_n_2303 = ({in2[3]} ^ {in1[27]});
 assign mul_34_17_n_2302 = ~({in2[7]} ^ {in1[10]});
 assign mul_34_17_n_2301 = ({in2[15]} ^ {in1[61]});
 assign mul_34_17_n_2300 = ({in2[11]} ^ {in1[22]});
 assign mul_34_17_n_2299 = ({in2[5]} ^ {in1[32]});
 assign mul_34_17_n_2298 = ~({in2[15]} ^ {in1[26]});
 assign mul_34_17_n_2297 = ~({in2[5]} ^ {in1[57]});
 assign mul_34_17_n_2296 = ~({in2[23]} ^ {in1[49]});
 assign mul_34_17_n_2294 = ~({in2[7]} ^ {in1[38]});
 assign mul_34_17_n_2293 = ~({in2[13]} ^ {in1[51]});
 assign mul_34_17_n_1694 = ~({in2[7]} ^ {in1[63]});
 assign mul_34_17_n_2291 = ({in2[7]} ^ {in1[15]});
 assign mul_34_17_n_2289 = ~({in2[3]} ^ {in1[18]});
 assign mul_34_17_n_2288 = ({in2[5]} ^ {in1[1]});
 assign mul_34_17_n_2286 = ~({in2[21]} ^ {in1[56]});
 assign mul_34_17_n_1693 = ~(mul_34_17_n_520 & mul_34_17_n_530);
 assign mul_34_17_n_2285 = ~({in2[17]} ^ {in1[29]});
 assign mul_34_17_n_2284 = ~({in2[19]} ^ {in1[57]});
 assign mul_34_17_n_2283 = ~({in2[5]} ^ {in1[40]});
 assign mul_34_17_n_2282 = ({in2[15]} ^ {in1[16]});
 assign mul_34_17_n_2280 = ~({in2[5]} ^ {in1[24]});
 assign mul_34_17_n_2279 = ({in2[17]} ^ {in1[15]});
 assign mul_34_17_n_2277 = ~({in2[13]} ^ {in1[53]});
 assign mul_34_17_n_2276 = ({in2[5]} ^ {in1[30]});
 assign mul_34_17_n_2275 = ({in2[15]} ^ {in1[18]});
 assign mul_34_17_n_2274 = ({in2[3]} ^ {in1[55]});
 assign mul_34_17_n_2273 = ({in2[3]} ^ {in1[30]});
 assign mul_34_17_n_2271 = ~({in2[7]} ^ {in1[34]});
 assign mul_34_17_n_2269 = ~({in2[13]} ^ {in1[2]});
 assign mul_34_17_n_2268 = ({in2[7]} ^ {in1[49]});
 assign mul_34_17_n_2267 = ~({in2[3]} ^ {in1[8]});
 assign mul_34_17_n_2265 = ~({in2[15]} ^ {in1[1]});
 assign mul_34_17_n_2264 = ~({in2[19]} ^ {in1[22]});
 assign mul_34_17_n_2263 = ~({in2[11]} ^ {in1[6]});
 assign mul_34_17_n_2262 = ~({in2[21]} ^ {in1[51]});
 assign mul_34_17_n_2261 = ({in2[25]} ^ {in1[29]});
 assign mul_34_17_n_2260 = ({in2[21]} ^ {in1[36]});
 assign mul_34_17_n_2259 = ({in2[21]} ^ {in1[10]});
 assign mul_34_17_n_2258 = ({in2[3]} ^ {in1[1]});
 assign mul_34_17_n_2256 = ~({in2[25]} ^ {in1[34]});
 assign mul_34_17_n_2255 = ({in2[23]} ^ {in1[34]});
 assign mul_34_17_n_2253 = ~({in2[7]} ^ {in1[52]});
 assign mul_34_17_n_2252 = ({in2[23]} ^ {in1[32]});
 assign mul_34_17_n_2250 = ~({in2[13]} ^ {in1[27]});
 assign mul_34_17_n_2248 = ~({in2[15]} ^ {in1[59]});
 assign mul_34_17_n_2247 = ({in2[7]} ^ {in1[46]});
 assign mul_34_17_n_2246 = ({in2[11]} ^ {in1[47]});
 assign mul_34_17_n_2245 = ({in2[13]} ^ {in1[7]});
 assign mul_34_17_n_2244 = ({in2[13]} ^ {in1[43]});
 assign mul_34_17_n_2242 = ~({in2[21]} ^ {in1[28]});
 assign mul_34_17_n_2241 = ~({in2[5]} ^ {in1[5]});
 assign mul_34_17_n_2240 = ({in2[15]} ^ {in1[60]});
 assign mul_34_17_n_2239 = ~(mul_34_17_n_517 & {in2[1]});
 assign mul_34_17_n_2238 = ({in2[15]} ^ {in1[19]});
 assign mul_34_17_n_2237 = ~({in2[7]} ^ {in1[53]});
 assign mul_34_17_n_2236 = ~({in2[17]} ^ {in1[57]});
 assign mul_34_17_n_2235 = ({in2[7]} ^ {in1[26]});
 assign mul_34_17_n_2234 = ~({in2[19]} ^ {in1[53]});
 assign mul_34_17_n_2232 = ~({in2[23]} ^ {in1[54]});
 assign mul_34_17_n_2231 = ~({in2[17]} ^ {in1[58]});
 assign mul_34_17_n_2230 = ~({in2[7]} ^ {in1[19]});
 assign mul_34_17_n_2229 = ~({in2[15]} ^ {in1[2]});
 assign mul_34_17_n_2228 = ({in2[3]} ^ {in1[29]});
 assign mul_34_17_n_2227 = ~({in2[5]} ^ {in1[17]});
 assign mul_34_17_n_2226 = ({in2[5]} ^ {in1[50]});
 assign mul_34_17_n_2224 = ~({in2[9]} ^ {in1[51]});
 assign mul_34_17_n_2223 = ({in2[13]} ^ {in1[20]});
 assign mul_34_17_n_2222 = ({in2[13]} ^ {in1[9]});
 assign mul_34_17_n_2221 = ({in2[13]} ^ {in1[19]});
 assign mul_34_17_n_2220 = ~({in2[9]} ^ {in1[8]});
 assign mul_34_17_n_2219 = ({in2[23]} ^ {in1[60]});
 assign mul_34_17_n_2218 = ({in2[19]} ^ {in1[1]});
 assign mul_34_17_n_2217 = ({in2[21]} ^ {in1[12]});
 assign mul_34_17_n_2216 = ~({in2[17]} ^ {in1[56]});
 assign mul_34_17_n_2215 = ~({in2[13]} ^ {in1[34]});
 assign mul_34_17_n_2214 = ~({in2[15]} ^ {in1[5]});
 assign mul_34_17_n_2213 = ({in2[9]} ^ {in1[24]});
 assign mul_34_17_n_2212 = ({in2[5]} ^ {in1[51]});
 assign mul_34_17_n_2211 = ({in2[23]} ^ {in1[17]});
 assign mul_34_17_n_2210 = ({in2[7]} ^ {in1[24]});
 assign mul_34_17_n_2209 = ({in2[11]} ^ {in1[52]});
 assign mul_34_17_n_2208 = ~({in2[13]} ^ {in1[60]});
 assign mul_34_17_n_2207 = ~({in2[13]} ^ {in1[62]});
 assign mul_34_17_n_2206 = ~({in2[13]} ^ {in1[61]});
 assign mul_34_17_n_2205 = ({in2[3]} ^ {in1[47]});
 assign mul_34_17_n_2204 = ~({in2[3]} ^ {in1[14]});
 assign mul_34_17_n_2203 = ({in2[11]} ^ {in1[26]});
 assign mul_34_17_n_2201 = ~({in2[21]} ^ {in1[62]});
 assign mul_34_17_n_2200 = ({in2[9]} ^ {in1[25]});
 assign mul_34_17_n_2199 = ~({in2[21]} ^ {in1[55]});
 assign mul_34_17_n_2197 = ~({in2[19]} ^ {in1[27]});
 assign mul_34_17_n_2196 = ({in2[7]} ^ {in1[14]});
 assign mul_34_17_n_2195 = ({in2[11]} ^ {in1[18]});
 assign mul_34_17_n_2194 = ~({in2[19]} ^ {in1[28]});
 assign mul_34_17_n_2193 = ({in2[17]} ^ {in1[20]});
 assign mul_34_17_n_2192 = ({in2[21]} ^ {in1[45]});
 assign mul_34_17_n_2191 = ~({in2[15]} ^ {in1[32]});
 assign mul_34_17_n_2190 = ({in2[17]} ^ {in1[18]});
 assign mul_34_17_n_2189 = ~({in2[5]} ^ {in1[56]});
 assign mul_34_17_n_2188 = ~({in2[11]} ^ {in1[10]});
 assign mul_34_17_n_2187 = ({in2[11]} ^ {in1[36]});
 assign mul_34_17_n_2186 = ~({in2[19]} ^ {in1[41]});
 assign mul_34_17_n_2185 = ({in2[3]} ^ {in1[19]});
 assign mul_34_17_n_1692 = ~(mul_34_17_n_525 | mul_34_17_n_529);
 assign mul_34_17_n_2184 = ~({in2[5]} ^ {in1[15]});
 assign mul_34_17_n_2183 = ~({in2[15]} ^ {in1[29]});
 assign mul_34_17_n_2181 = ~({in2[13]} ^ {in1[6]});
 assign mul_34_17_n_2179 = ~({in2[9]} ^ {in1[31]});
 assign mul_34_17_n_2178 = ~({in2[13]} ^ {in1[58]});
 assign mul_34_17_n_2176 = ~({in2[3]} ^ {in1[58]});
 assign mul_34_17_n_2175 = ({in2[3]} ^ {in1[39]});
 assign mul_34_17_n_2174 = ({in2[5]} ^ {in1[10]});
 assign mul_34_17_n_2173 = ~({in2[19]} ^ {in1[20]});
 assign mul_34_17_n_2172 = ~({in2[21]} ^ {in1[23]});
 assign mul_34_17_n_2171 = ~({in2[19]} ^ {in1[19]});
 assign mul_34_17_n_2170 = ({in2[23]} ^ {in1[5]});
 assign mul_34_17_n_2168 = ~({in2[5]} ^ {in1[54]});
 assign mul_34_17_n_2167 = ~({in2[19]} ^ {in1[3]});
 assign mul_34_17_n_2166 = ~({in2[15]} ^ {in1[3]});
 assign mul_34_17_n_2164 = ~({in2[3]} ^ {in1[38]});
 assign mul_34_17_n_2163 = ({in2[25]} ^ {in1[28]});
 assign mul_34_17_n_2161 = ~({in2[3]} ^ {in1[9]});
 assign mul_34_17_n_2160 = ~({in2[15]} ^ {in1[4]});
 assign mul_34_17_n_2159 = ({in2[11]} ^ {in1[53]});
 assign mul_34_17_n_1691 = ({in2[3]} ^ {in1[63]});
 assign mul_34_17_n_2157 = ({in2[17]} ^ {in1[21]});
 assign mul_34_17_n_2156 = ~({in2[21]} ^ {in1[4]});
 assign mul_34_17_n_2155 = ~({in2[15]} ^ {in1[53]});
 assign mul_34_17_n_2154 = ~({in2[23]} ^ {in1[37]});
 assign mul_34_17_n_2152 = ~({in2[5]} ^ {in1[42]});
 assign mul_34_17_n_2151 = ({in2[17]} ^ {in1[38]});
 assign mul_34_17_n_2150 = ~({in2[19]} ^ {in1[7]});
 assign mul_34_17_n_2149 = ({in2[3]} ^ {in1[10]});
 assign mul_34_17_n_2148 = ({in2[23]} ^ {in1[56]});
 assign mul_34_17_n_2147 = ~({in2[5]} ^ {in1[36]});
 assign mul_34_17_n_2146 = ({in2[21]} ^ {in1[31]});
 assign mul_34_17_n_2145 = ({in2[23]} ^ {in1[9]});
 assign mul_34_17_n_2144 = ~({in2[17]} ^ {in1[8]});
 assign mul_34_17_n_2142 = ~({in2[7]} ^ {in1[59]});
 assign mul_34_17_n_2141 = ({in2[17]} ^ {in1[39]});
 assign mul_34_17_n_2139 = ~({in2[17]} ^ {in1[30]});
 assign mul_34_17_n_2138 = ({in2[3]} ^ {in1[61]});
 assign mul_34_17_n_2136 = ~({in2[21]} ^ {in1[60]});
 assign mul_34_17_n_2135 = ({in2[3]} ^ {in1[45]});
 assign mul_34_17_n_2134 = ({in2[9]} ^ {in1[47]});
 assign mul_34_17_n_2133 = ({in2[23]} ^ {in1[14]});
 assign mul_34_17_n_2132 = ~({in2[7]} ^ {in1[9]});
 assign mul_34_17_n_2131 = ({in2[19]} ^ {in1[49]});
 assign mul_34_17_n_2130 = ({in2[11]} ^ {in1[21]});
 assign mul_34_17_n_2129 = ~({in2[9]} ^ {in1[40]});
 assign mul_34_17_n_2127 = ({in2[19]} ^ {in1[31]});
 assign mul_34_17_n_2125 = ~({in2[11]} ^ {in1[15]});
 assign mul_34_17_n_2124 = ({in2[3]} ^ {in1[4]});
 assign mul_34_17_n_2123 = ({in2[11]} ^ {in1[51]});
 assign mul_34_17_n_2121 = ~({in2[7]} ^ {in1[4]});
 assign mul_34_17_n_2120 = ({in2[17]} ^ {in1[16]});
 assign mul_34_17_n_2119 = ({in2[3]} ^ {in1[49]});
 assign mul_34_17_n_2118 = ({in2[15]} ^ {in1[17]});
 assign mul_34_17_n_2116 = ({in2[5]} ^ {in1[28]});
 assign mul_34_17_n_2115 = ({in2[3]} ^ {in1[51]});
 assign mul_34_17_n_2114 = ({in2[21]} ^ {in1[40]});
 assign mul_34_17_n_2112 = ~({in2[11]} ^ {in1[49]});
 assign mul_34_17_n_2111 = ~({in2[7]} ^ {in1[55]});
 assign mul_34_17_n_2110 = ~({in2[11]} ^ {in1[9]});
 assign mul_34_17_n_2109 = ({in2[15]} ^ {in1[24]});
 assign mul_34_17_n_2108 = ({in2[5]} ^ {in1[26]});
 assign mul_34_17_n_2107 = ~({in2[21]} ^ {in1[50]});
 assign mul_34_17_n_2105 = ~({in2[11]} ^ {in1[57]});
 assign mul_34_17_n_2103 = ~({in2[3]} ^ {in1[6]});
 assign mul_34_17_n_2102 = ~({in2[15]} ^ {in1[57]});
 assign mul_34_17_n_2101 = ({in2[7]} ^ {in1[32]});
 assign mul_34_17_n_2100 = ({in2[5]} ^ {in1[7]});
 assign mul_34_17_n_2099 = ~({in2[17]} ^ {in1[28]});
 assign mul_34_17_n_2098 = ~({in2[11]} ^ {in1[38]});
 assign mul_34_17_n_2096 = ~({in2[25]} ^ {in1[55]});
 assign mul_34_17_n_2095 = ({in2[3]} ^ {in1[56]});
 assign mul_34_17_n_2093 = ~({in2[17]} ^ {in1[32]});
 assign mul_34_17_n_2091 = ~({in2[21]} ^ {in1[27]});
 assign mul_34_17_n_2090 = ~({in2[23]} ^ {in1[47]});
 assign mul_34_17_n_2089 = ~({in2[9]} ^ {in1[16]});
 assign mul_34_17_n_2088 = ({in2[23]} ^ {in1[8]});
 assign mul_34_17_n_2087 = ~({in2[5]} ^ {in1[19]});
 assign mul_34_17_n_2085 = ~({in2[9]} ^ {in1[3]});
 assign mul_34_17_n_2084 = ~({in2[7]} ^ {in1[11]});
 assign mul_34_17_n_2083 = ~({in2[23]} ^ {in1[39]});
 assign mul_34_17_n_2082 = ({in2[19]} ^ {in1[36]});
 assign mul_34_17_n_2080 = ({in2[5]} ^ {in1[3]});
 assign mul_34_17_n_2079 = ~({in2[17]} ^ {in1[60]});
 assign mul_34_17_n_2077 = ({in2[23]} ^ {in1[16]});
 assign mul_34_17_n_2076 = ~({in2[7]} ^ {in1[37]});
 assign mul_34_17_n_2074 = ({in2[19]} ^ {in1[2]});
 assign mul_34_17_n_2072 = ({in2[3]} ^ {in1[40]});
 assign mul_34_17_n_2071 = ({in2[19]} ^ {in1[39]});
 assign mul_34_17_n_2070 = ({in2[19]} ^ {in1[37]});
 assign mul_34_17_n_2068 = ~({in2[21]} ^ {in1[22]});
 assign mul_34_17_n_2067 = ~({in2[9]} ^ {in1[62]});
 assign mul_34_17_n_2066 = ~({in2[13]} ^ {in1[29]});
 assign mul_34_17_n_2064 = ({in2[9]} ^ {in1[53]});
 assign mul_34_17_n_2063 = ({in2[9]} ^ {in1[52]});
 assign mul_34_17_n_2061 = ~({in2[19]} ^ {in1[58]});
 assign mul_34_17_n_2060 = ~({in2[19]} ^ {in1[25]});
 assign mul_34_17_n_2059 = ({in2[23]} ^ {in1[57]});
 assign mul_34_17_n_2058 = ~({in2[15]} ^ {in1[13]});
 assign mul_34_17_n_2057 = ~({in2[17]} ^ {in1[54]});
 assign mul_34_17_n_2056 = ({in2[13]} ^ {in1[17]});
 assign mul_34_17_n_2055 = ~({in2[23]} ^ {in1[21]});
 assign mul_34_17_n_2054 = ({in2[9]} ^ {in1[49]});
 assign mul_34_17_n_2053 = ~({in2[11]} ^ {in1[33]});
 assign mul_34_17_n_2052 = ~({in2[11]} ^ {in1[32]});
 assign mul_34_17_n_2050 = ({in2[9]} ^ {in1[41]});
 assign mul_34_17_n_2049 = ~({in2[19]} ^ {in1[52]});
 assign mul_34_17_n_2048 = ~({in2[17]} ^ {in1[6]});
 assign mul_34_17_n_2047 = ({in2[9]} ^ {in1[33]});
 assign mul_34_17_n_2045 = ~({in2[11]} ^ {in1[39]});
 assign mul_34_17_n_2044 = ({in2[7]} ^ {in1[43]});
 assign mul_34_17_n_2043 = ({in2[9]} ^ {in1[4]});
 assign mul_34_17_n_2042 = ~({in2[21]} ^ {in1[52]});
 assign mul_34_17_n_2040 = ~({in2[23]} ^ {in1[43]});
 assign mul_34_17_n_2039 = ({in2[7]} ^ {in1[35]});
 assign mul_34_17_n_2038 = ~({in2[17]} ^ {in1[25]});
 assign mul_34_17_n_2037 = ~({in2[13]} ^ {in1[37]});
 assign mul_34_17_n_2036 = ({in2[9]} ^ {in1[30]});
 assign mul_34_17_n_2034 = ~({in2[3]} ^ {in1[16]});
 assign mul_34_17_n_2032 = ~({in2[9]} ^ {in1[29]});
 assign mul_34_17_n_2031 = ~({in2[19]} ^ {in1[51]});
 assign mul_34_17_n_2030 = ~({in2[17]} ^ {in1[23]});
 assign mul_34_17_n_2029 = ~({in2[7]} ^ {in1[16]});
 assign mul_34_17_n_2028 = ({in2[5]} ^ {in1[8]});
 assign mul_34_17_n_1690 = ~(mul_34_17_n_519 & mul_34_17_n_521);
 assign mul_34_17_n_2026 = ~({in2[23]} ^ {in1[36]});
 assign mul_34_17_n_2024 = ({in2[3]} ^ {in1[20]});
 assign mul_34_17_n_2022 = ~({in2[21]} ^ {in1[42]});
 assign mul_34_17_n_2020 = ~({in2[21]} ^ {in1[29]});
 assign mul_34_17_n_2019 = ~({in2[9]} ^ {in1[14]});
 assign mul_34_17_n_2018 = ({in2[3]} ^ {in1[32]});
 assign mul_34_17_n_2016 = ({in2[3]} ^ {in1[60]});
 assign mul_34_17_n_2015 = ~({in2[3]} ^ {in1[21]});
 assign mul_34_17_n_2013 = ~({in2[23]} ^ {in1[18]});
 assign mul_34_17_n_2012 = ~({in2[21]} ^ {in1[18]});
 assign mul_34_17_n_2011 = ({in2[7]} ^ {in1[25]});
 assign mul_34_17_n_2009 = ~({in2[19]} ^ {in1[46]});
 assign mul_34_17_n_2008 = ({in2[21]} ^ {in1[37]});
 assign mul_34_17_n_2007 = ({in2[5]} ^ {in1[33]});
 assign mul_34_17_n_2006 = ~({in2[7]} ^ {in1[21]});
 assign mul_34_17_n_2005 = ~({in2[23]} ^ {in1[19]});
 assign mul_34_17_n_2004 = ~({in2[5]} ^ {in1[18]});
 assign mul_34_17_n_2003 = ~({in2[5]} ^ {in1[38]});
 assign mul_34_17_n_2001 = ~({in2[13]} ^ {in1[15]});
 assign mul_34_17_n_1999 = ~({in2[23]} ^ {in1[28]});
 assign mul_34_17_n_1998 = ~({in2[21]} ^ {in1[53]});
 assign mul_34_17_n_1997 = ~({in2[19]} ^ {in1[9]});
 assign mul_34_17_n_1996 = ~({in2[11]} ^ {in1[5]});
 assign mul_34_17_n_1995 = ({in2[21]} ^ {in1[59]});
 assign mul_34_17_n_1994 = ({in2[7]} ^ {in1[13]});
 assign mul_34_17_n_1993 = ({in2[21]} ^ {in1[33]});
 assign mul_34_17_n_1992 = ({in2[7]} ^ {in1[7]});
 assign mul_34_17_n_1991 = ~({in2[9]} ^ {in1[56]});
 assign mul_34_17_n_1990 = ({in2[5]} ^ {in1[49]});
 assign mul_34_17_n_1989 = ({in2[17]} ^ {in1[51]});
 assign mul_34_17_n_1988 = ~({in2[15]} ^ {in1[27]});
 assign mul_34_17_n_1986 = ~({in2[9]} ^ {in1[34]});
 assign mul_34_17_n_1984 = ({in2[17]} ^ {in1[5]});
 assign mul_34_17_n_1983 = ~({in2[21]} ^ {in1[19]});
 assign mul_34_17_n_1981 = ~({in2[23]} ^ {in1[45]});
 assign mul_34_17_n_1979 = ~({in2[13]} ^ {in1[33]});
 assign mul_34_17_n_1978 = ({in2[21]} ^ {in1[46]});
 assign mul_34_17_n_1976 = ~({in2[13]} ^ {in1[55]});
 assign mul_34_17_n_1974 = ~({in2[25]} ^ {in1[12]});
 assign mul_34_17_n_1973 = ({in2[17]} ^ {in1[14]});
 assign mul_34_17_n_1972 = ({in2[11]} ^ {in1[29]});
 assign mul_34_17_n_1971 = ({in2[11]} ^ {in1[27]});
 assign mul_34_17_n_1969 = ~({in2[21]} ^ {in1[8]});
 assign mul_34_17_n_1968 = ({in2[3]} ^ {in1[35]});
 assign mul_34_17_n_1967 = ~({in2[23]} ^ {in1[48]});
 assign mul_34_17_n_1965 = ~({in2[15]} ^ {in1[45]});
 assign mul_34_17_n_1963 = ~({in2[9]} ^ {in1[20]});
 assign mul_34_17_n_1962 = ({in2[13]} ^ {in1[25]});
 assign mul_34_17_n_1961 = ~({in2[15]} ^ {in1[30]});
 assign mul_34_17_n_1960 = ({in2[9]} ^ {in1[46]});
 assign mul_34_17_n_1958 = ~({in2[25]} ^ {in1[16]});
 assign mul_34_17_n_1957 = ({in2[11]} ^ {in1[42]});
 assign mul_34_17_n_1956 = ({in2[15]} ^ {in1[21]});
 assign mul_34_17_n_1955 = ({in2[11]} ^ {in1[43]});
 assign mul_34_17_n_1954 = ~({in2[9]} ^ {in1[39]});
 assign mul_34_17_n_1952 = ~({in2[17]} ^ {in1[46]});
 assign mul_34_17_n_1950 = ~({in2[23]} ^ {in1[22]});
 assign mul_34_17_n_1948 = ({in2[11]} ^ {in1[37]});
 assign mul_34_17_n_1947 = ({in2[17]} ^ {in1[37]});
 assign mul_34_17_n_1946 = ~({in2[5]} ^ {in1[37]});
 assign mul_34_17_n_1945 = ({in2[5]} ^ {in1[60]});
 assign mul_34_17_n_1944 = ~({in2[21]} ^ {in1[7]});
 assign mul_34_17_n_1943 = ~({in2[15]} ^ {in1[54]});
 assign mul_34_17_n_1941 = ~({in2[19]} ^ {in1[50]});
 assign mul_34_17_n_1940 = ~({in2[13]} ^ {in1[56]});
 assign mul_34_17_n_1938 = ~({in2[17]} ^ {in1[45]});
 assign mul_34_17_n_1937 = ~({in2[23]} ^ {in1[25]});
 assign mul_34_17_n_1935 = ~({in2[5]} ^ {in1[27]});
 assign mul_34_17_n_1934 = ({in2[11]} ^ {in1[25]});
 assign mul_34_17_n_1933 = ~({in2[17]} ^ {in1[24]});
 assign mul_34_17_n_1932 = ~({in2[13]} ^ {in1[35]});
 assign mul_34_17_n_1931 = ({in2[5]} ^ {in1[31]});
 assign mul_34_17_n_1930 = ({in2[7]} ^ {in1[41]});
 assign mul_34_17_n_1929 = ~({in2[21]} ^ {in1[54]});
 assign mul_34_17_n_1928 = ({in2[7]} ^ {in1[30]});
 assign mul_34_17_n_1927 = ~({in2[11]} ^ {in1[31]});
 assign mul_34_17_n_1926 = ({in2[19]} ^ {in1[59]});
 assign mul_34_17_n_1925 = ({in2[7]} ^ {in1[29]});
 assign mul_34_17_n_1923 = ~({in2[17]} ^ {in1[52]});
 assign mul_34_17_n_1922 = ~({in2[19]} ^ {in1[56]});
 assign mul_34_17_n_1921 = ~({in2[23]} ^ {in1[20]});
 assign mul_34_17_n_1919 = ~({in2[3]} ^ {in1[34]});
 assign mul_34_17_n_1918 = ~({in2[19]} ^ {in1[5]});
 assign mul_34_17_n_1917 = ~({in2[3]} ^ {in1[13]});
 assign mul_34_17_n_1916 = ~({in2[23]} ^ {in1[40]});
 assign mul_34_17_n_1914 = ({in2[21]} ^ {in1[2]});
 assign mul_34_17_n_1913 = ~({in2[17]} ^ {in1[61]});
 assign mul_34_17_n_1912 = ~({in2[19]} ^ {in1[29]});
 assign mul_34_17_n_1911 = ~({in2[11]} ^ {in1[13]});
 assign mul_34_17_n_1910 = ~({in2[11]} ^ {in1[12]});
 assign mul_34_17_n_1909 = ~({in2[19]} ^ {in1[4]});
 assign mul_34_17_n_1908 = ({in2[17]} ^ {in1[10]});
 assign mul_34_17_n_1907 = ~({in2[9]} ^ {in1[60]});
 assign mul_34_17_n_1906 = ~({in2[23]} ^ {in1[38]});
 assign mul_34_17_n_1904 = ~({in2[7]} ^ {in1[36]});
 assign mul_34_17_n_1903 = ({in2[15]} ^ {in1[49]});
 assign mul_34_17_n_1902 = ~({in2[17]} ^ {in1[26]});
 assign mul_34_17_n_1689 = ({in2[15]} ^ {in1[63]});
 assign mul_34_17_n_1900 = ({in2[13]} ^ {in1[50]});
 assign mul_34_17_n_1898 = ~({in2[7]} ^ {in1[56]});
 assign mul_34_17_n_1896 = ~({in2[13]} ^ {in1[41]});
 assign mul_34_17_n_1895 = ~({in2[17]} ^ {in1[7]});
 assign mul_34_17_n_1894 = ~({in2[19]} ^ {in1[10]});
 assign mul_34_17_n_1893 = ~({in2[5]} ^ {in1[20]});
 assign mul_34_17_n_1892 = ~({in2[19]} ^ {in1[44]});
 assign mul_34_17_n_1891 = ~({in2[13]} ^ {in1[12]});
 assign mul_34_17_n_1890 = ({in2[7]} ^ {in1[44]});
 assign mul_34_17_n_1889 = ({in2[23]} ^ {in1[4]});
 assign mul_34_17_n_1887 = ~({in2[13]} ^ {in1[32]});
 assign mul_34_17_n_1886 = ({in2[5]} ^ {in1[44]});
 assign mul_34_17_n_1884 = ~({in2[23]} ^ {in1[51]});
 assign mul_34_17_n_1883 = ~({in2[7]} ^ {in1[18]});
 assign mul_34_17_n_1881 = ~({in2[23]} ^ {in1[2]});
 assign mul_34_17_n_1879 = ~({in2[15]} ^ {in1[10]});
 assign mul_34_17_n_1878 = ({in2[5]} ^ {in1[52]});
 assign mul_34_17_n_1877 = ({in2[21]} ^ {in1[15]});
 assign mul_34_17_n_1876 = ({in2[15]} ^ {in1[51]});
 assign mul_34_17_n_1875 = ({in2[3]} ^ {in1[36]});
 assign mul_34_17_n_1874 = ~({in2[21]} ^ {in1[5]});
 assign mul_34_17_n_1873 = ({in2[21]} ^ {in1[21]});
 assign mul_34_17_n_1872 = ~({in2[3]} ^ {in1[22]});
 assign mul_34_17_n_1871 = ({in2[15]} ^ {in1[40]});
 assign mul_34_17_n_1870 = ({in2[5]} ^ {in1[43]});
 assign mul_34_17_n_1869 = ~({in2[7]} ^ {in1[3]});
 assign mul_34_17_n_1867 = ~({in2[17]} ^ {in1[33]});
 assign mul_34_17_n_1866 = ({in2[13]} ^ {in1[24]});
 assign mul_34_17_n_1864 = ~({in2[5]} ^ {in1[6]});
 assign mul_34_17_n_1863 = ({in2[15]} ^ {in1[15]});
 assign mul_34_17_n_1861 = ~({in2[7]} ^ {in1[23]});
 assign mul_34_17_n_1860 = ({in2[11]} ^ {in1[41]});
 assign mul_34_17_n_1859 = ~({in2[17]} ^ {in1[22]});
 assign mul_34_17_n_1858 = ({in2[23]} ^ {in1[3]});
 assign mul_34_17_n_1857 = ~({in2[9]} ^ {in1[17]});
 assign mul_34_17_n_1856 = ~({in2[11]} ^ {in1[11]});
 assign mul_34_17_n_1855 = ~({in2[9]} ^ {in1[55]});
 assign mul_34_17_n_1854 = ~({in2[11]} ^ {in1[8]});
 assign mul_34_17_n_1853 = ({in2[17]} ^ {in1[11]});
 assign mul_34_17_n_1852 = ~({in2[19]} ^ {in1[8]});
 assign mul_34_17_n_1851 = ~({in2[15]} ^ {in1[58]});
 assign mul_34_17_n_1850 = ({in2[7]} ^ {in1[48]});
 assign mul_34_17_n_1849 = ({in2[23]} ^ {in1[33]});
 assign mul_34_17_n_1848 = ({in2[7]} ^ {in1[45]});
 assign mul_34_17_n_1847 = ({in2[11]} ^ {in1[16]});
 assign mul_34_17_n_1846 = ({in2[7]} ^ {in1[1]});
 assign mul_34_17_n_1844 = ~({in2[23]} ^ {in1[59]});
 assign mul_34_17_n_1842 = ~({in2[23]} ^ {in1[58]});
 assign mul_34_17_n_1841 = ({in2[11]} ^ {in1[2]});
 assign mul_34_17_n_1840 = ({in2[21]} ^ {in1[34]});
 assign mul_34_17_n_1839 = ({in2[1]} ^ {in1[5]});
 assign mul_34_17_n_1838 = ({in2[1]} ^ {in1[43]});
 assign mul_34_17_n_1837 = ({in2[1]} ^ {in1[10]});
 assign mul_34_17_n_1836 = ({in2[1]} ^ {in1[44]});
 assign mul_34_17_n_1835 = ({in2[1]} ^ {in1[11]});
 assign mul_34_17_n_1834 = ({in2[1]} ^ {in1[38]});
 assign mul_34_17_n_1833 = ({in2[1]} ^ {in1[24]});
 assign mul_34_17_n_1832 = ({in2[1]} ^ {in1[23]});
 assign mul_34_17_n_1831 = ({in2[25]} ^ {in1[9]});
 assign mul_34_17_n_1830 = ({in2[1]} ^ {in1[34]});
 assign mul_34_17_n_1829 = ({in2[1]} ^ {in1[40]});
 assign mul_34_17_n_1828 = ({in2[1]} ^ {in1[25]});
 assign mul_34_17_n_1827 = ({in2[1]} ^ {in1[42]});
 assign mul_34_17_n_1826 = ({in2[1]} ^ {in1[52]});
 assign mul_34_17_n_1825 = ({in2[1]} ^ {in1[29]});
 assign mul_34_17_n_1824 = ({in2[1]} ^ {in1[1]});
 assign mul_34_17_n_1823 = ({in2[1]} ^ {in1[54]});
 assign mul_34_17_n_1822 = ({in2[1]} ^ {in1[51]});
 assign mul_34_17_n_1821 = ({in2[1]} ^ {in1[30]});
 assign mul_34_17_n_1820 = ({in2[1]} ^ {in1[26]});
 assign mul_34_17_n_1819 = ({in2[1]} ^ {in1[4]});
 assign mul_34_17_n_1818 = ({in2[1]} ^ {in1[27]});
 assign mul_34_17_n_1817 = ({in2[1]} ^ {in1[7]});
 assign mul_34_17_n_1816 = ({in2[1]} ^ {in1[53]});
 assign mul_34_17_n_1815 = ({in2[1]} ^ {in1[8]});
 assign mul_34_17_n_1814 = ({in2[1]} ^ {in1[59]});
 assign mul_34_17_n_1813 = ({in2[1]} ^ {in1[36]});
 assign mul_34_17_n_1812 = ({in2[1]} ^ {in1[46]});
 assign mul_34_17_n_1811 = ({in2[1]} ^ {in1[28]});
 assign mul_34_17_n_1810 = ({in2[1]} ^ {in1[2]});
 assign mul_34_17_n_1809 = ({in2[1]} ^ {in1[15]});
 assign mul_34_17_n_1808 = ({in2[1]} ^ {in1[9]});
 assign mul_34_17_n_1807 = ({in2[1]} ^ {in1[20]});
 assign mul_34_17_n_1806 = ({in2[1]} ^ {in1[50]});
 assign mul_34_17_n_1805 = ({in2[1]} ^ {in1[12]});
 assign mul_34_17_n_1804 = ({in2[1]} ^ {in1[17]});
 assign mul_34_17_n_1803 = ({in2[1]} ^ {in1[13]});
 assign mul_34_17_n_1802 = ({in2[1]} ^ {in1[31]});
 assign mul_34_17_n_1801 = ({in2[1]} ^ {in1[16]});
 assign mul_34_17_n_1800 = ({in2[1]} ^ {in1[14]});
 assign mul_34_17_n_1799 = ({in2[1]} ^ {in1[48]});
 assign mul_34_17_n_1798 = ({in2[1]} ^ {in1[19]});
 assign mul_34_17_n_1797 = ({in2[1]} ^ {in1[37]});
 assign mul_34_17_n_1796 = ({in2[1]} ^ {in1[18]});
 assign mul_34_17_n_1795 = ({in2[1]} ^ {in1[62]});
 assign mul_34_17_n_1794 = ({in2[1]} ^ {in1[35]});
 assign mul_34_17_n_1793 = ({in2[1]} ^ {in1[6]});
 assign mul_34_17_n_1792 = ({in2[1]} ^ {in1[41]});
 assign mul_34_17_n_1791 = ({in2[1]} ^ {in1[60]});
 assign mul_34_17_n_1790 = ({in2[1]} ^ {in1[56]});
 assign mul_34_17_n_1789 = ({in2[1]} ^ {in1[61]});
 assign mul_34_17_n_1788 = ({in2[1]} ^ {in1[39]});
 assign mul_34_17_n_1787 = ({in2[1]} ^ {in1[55]});
 assign mul_34_17_n_1786 = ({in2[1]} ^ {in1[45]});
 assign mul_34_17_n_1785 = ({in2[1]} ^ {in1[32]});
 assign mul_34_17_n_1784 = ({in2[1]} ^ {in1[3]});
 assign mul_34_17_n_1688 = ({in2[1]} ^ {in1[63]});
 assign mul_34_17_n_1783 = ({in2[1]} ^ {in1[47]});
 assign mul_34_17_n_1782 = ({in2[1]} ^ {in1[21]});
 assign mul_34_17_n_1781 = ({in2[1]} ^ {in1[22]});
 assign mul_34_17_n_1780 = ({in2[1]} ^ {in1[49]});
 assign mul_34_17_n_1779 = ({in2[1]} ^ {in1[33]});
 assign mul_34_17_n_1778 = ({in2[1]} ^ {in1[58]});
 assign mul_34_17_n_1777 = ({in2[1]} ^ {in1[57]});
 assign mul_34_17_n_1776 = ({in2[25]} ^ {in1[59]});
 assign mul_34_17_n_1775 = ~({in2[25]} ^ {in1[25]});
 assign mul_34_17_n_1774 = ({in2[25]} ^ {in1[14]});
 assign mul_34_17_n_1772 = ~({in2[25]} ^ {in1[37]});
 assign mul_34_17_n_1771 = ({in2[25]} ^ {in1[32]});
 assign mul_34_17_n_1770 = ~({in2[25]} ^ {in1[23]});
 assign mul_34_17_n_1768 = ~({in2[25]} ^ {in1[4]});
 assign mul_34_17_n_1766 = ~({in2[25]} ^ {in1[54]});
 assign mul_34_17_n_1765 = ({in2[25]} ^ {in1[31]});
 assign mul_34_17_n_1764 = ({in2[25]} ^ {in1[33]});
 assign mul_34_17_n_1763 = ({in2[25]} ^ {in1[58]});
 assign mul_34_17_n_1761 = ({in2[25]} ^ {in1[26]});
 assign mul_34_17_n_1760 = ({in2[25]} ^ {in1[53]});
 assign mul_34_17_n_1759 = ({in2[25]} ^ {in1[10]});
 assign mul_34_17_n_1758 = ~({in2[25]} ^ {in1[19]});
 assign mul_34_17_n_1757 = ({in2[23]} ^ {in2[24]});
 assign mul_34_17_n_1755 = ({in2[21]} ^ {in2[22]});
 assign mul_34_17_n_1753 = ({in2[19]} ^ {in2[20]});
 assign mul_34_17_n_1751 = ({in2[7]} ^ {in2[8]});
 assign mul_34_17_n_1749 = ({in2[5]} ^ {in2[6]});
 assign mul_34_17_n_1747 = ({in2[3]} ^ {in2[4]});
 assign mul_34_17_n_1745 = ({in2[1]} ^ {in2[2]});
 assign mul_34_17_n_1743 = ({in2[13]} ^ {in2[14]});
 assign mul_34_17_n_1741 = ({in2[15]} ^ {in2[16]});
 assign mul_34_17_n_1739 = ({in2[9]} ^ {in2[10]});
 assign mul_34_17_n_1737 = ({in2[11]} ^ {in2[12]});
 assign mul_34_17_n_1735 = ({in2[17]} ^ {in2[18]});
 assign mul_34_17_n_1685 = ~mul_34_17_n_1684;
 assign mul_34_17_n_1682 = ~mul_34_17_n_1681;
 assign mul_34_17_n_1679 = ~mul_34_17_n_1678;
 assign mul_34_17_n_1676 = ~mul_34_17_n_1675;
 assign mul_34_17_n_1674 = ~mul_34_17_n_1673;
 assign mul_34_17_n_1672 = ~mul_34_17_n_1671;
 assign mul_34_17_n_1668 = ~mul_34_17_n_1667;
 assign mul_34_17_n_1666 = ~mul_34_17_n_1665;
 assign mul_34_17_n_1658 = ~mul_34_17_n_1657;
 assign mul_34_17_n_1656 = ~mul_34_17_n_1655;
 assign mul_34_17_n_1653 = ~mul_34_17_n_1652;
 assign mul_34_17_n_1650 = ~mul_34_17_n_1649;
 assign mul_34_17_n_1641 = ~mul_34_17_n_1640;
 assign mul_34_17_n_1637 = ~mul_34_17_n_1636;
 assign mul_34_17_n_1635 = ~mul_34_17_n_1634;
 assign mul_34_17_n_1625 = ~mul_34_17_n_1624;
 assign mul_34_17_n_1621 = ~mul_34_17_n_1620;
 assign mul_34_17_n_1618 = ~mul_34_17_n_1617;
 assign mul_34_17_n_1613 = ~mul_34_17_n_1612;
 assign mul_34_17_n_1610 = ~mul_34_17_n_1609;
 assign mul_34_17_n_1608 = ~mul_34_17_n_1607;
 assign mul_34_17_n_1604 = ~mul_34_17_n_1603;
 assign mul_34_17_n_1602 = ~mul_34_17_n_1601;
 assign mul_34_17_n_1588 = ~mul_34_17_n_1587;
 assign mul_34_17_n_1582 = ~mul_34_17_n_1581;
 assign mul_34_17_n_1580 = ~mul_34_17_n_1579;
 assign mul_34_17_n_1564 = ~mul_34_17_n_1563;
 assign mul_34_17_n_1557 = ~mul_34_17_n_1556;
 assign mul_34_17_n_1554 = ~mul_34_17_n_1553;
 assign mul_34_17_n_1552 = ~mul_34_17_n_1551;
 assign mul_34_17_n_1547 = ~mul_34_17_n_1546;
 assign mul_34_17_n_1540 = ~mul_34_17_n_1539;
 assign mul_34_17_n_1538 = ~mul_34_17_n_1537;
 assign mul_34_17_n_1533 = ~mul_34_17_n_1532;
 assign mul_34_17_n_1528 = ~mul_34_17_n_1527;
 assign mul_34_17_n_1518 = ~mul_34_17_n_1517;
 assign mul_34_17_n_1516 = ~mul_34_17_n_1515;
 assign mul_34_17_n_1511 = ~mul_34_17_n_1510;
 assign mul_34_17_n_1508 = ~mul_34_17_n_1507;
 assign mul_34_17_n_1504 = ~mul_34_17_n_1503;
 assign mul_34_17_n_1502 = ~mul_34_17_n_1501;
 assign mul_34_17_n_1499 = ~mul_34_17_n_1498;
 assign mul_34_17_n_1494 = ~mul_34_17_n_1493;
 assign mul_34_17_n_1492 = ~mul_34_17_n_1491;
 assign mul_34_17_n_1490 = ~mul_34_17_n_1489;
 assign mul_34_17_n_1487 = ~mul_34_17_n_1486;
 assign mul_34_17_n_1484 = ~mul_34_17_n_1483;
 assign mul_34_17_n_1475 = ~mul_34_17_n_1474;
 assign mul_34_17_n_1470 = ~mul_34_17_n_1469;
 assign mul_34_17_n_1465 = ~mul_34_17_n_1464;
 assign mul_34_17_n_1462 = ~mul_34_17_n_1461;
 assign mul_34_17_n_1455 = ~mul_34_17_n_1454;
 assign mul_34_17_n_1447 = ~mul_34_17_n_1446;
 assign mul_34_17_n_1445 = ~mul_34_17_n_1444;
 assign mul_34_17_n_1440 = ~mul_34_17_n_1439;
 assign mul_34_17_n_1433 = ~mul_34_17_n_1432;
 assign mul_34_17_n_1431 = ~mul_34_17_n_1430;
 assign mul_34_17_n_1425 = ~mul_34_17_n_1424;
 assign mul_34_17_n_1421 = ~mul_34_17_n_1420;
 assign mul_34_17_n_1418 = ~mul_34_17_n_1417;
 assign mul_34_17_n_1416 = ~mul_34_17_n_1415;
 assign mul_34_17_n_1408 = ~mul_34_17_n_1407;
 assign mul_34_17_n_1406 = ~mul_34_17_n_1405;
 assign mul_34_17_n_1404 = ~mul_34_17_n_1403;
 assign mul_34_17_n_1402 = ~mul_34_17_n_1401;
 assign mul_34_17_n_1400 = ~mul_34_17_n_1399;
 assign mul_34_17_n_1394 = ~mul_34_17_n_1393;
 assign mul_34_17_n_1388 = ~mul_34_17_n_1387;
 assign mul_34_17_n_1383 = ~mul_34_17_n_1382;
 assign mul_34_17_n_1380 = ~mul_34_17_n_1379;
 assign mul_34_17_n_1377 = ~mul_34_17_n_1376;
 assign mul_34_17_n_1371 = ~mul_34_17_n_1370;
 assign mul_34_17_n_1365 = ~mul_34_17_n_1364;
 assign mul_34_17_n_1361 = ~mul_34_17_n_1360;
 assign mul_34_17_n_1359 = ~mul_34_17_n_1358;
 assign mul_34_17_n_1346 = ~mul_34_17_n_1345;
 assign mul_34_17_n_1339 = ~mul_34_17_n_1338;
 assign mul_34_17_n_1336 = ~mul_34_17_n_1335;
 assign mul_34_17_n_1334 = ~mul_34_17_n_1333;
 assign mul_34_17_n_1324 = ~mul_34_17_n_1323;
 assign mul_34_17_n_1320 = ~mul_34_17_n_1319;
 assign mul_34_17_n_1318 = ~mul_34_17_n_1317;
 assign mul_34_17_n_1315 = ~mul_34_17_n_1314;
 assign mul_34_17_n_1313 = ~mul_34_17_n_1312;
 assign mul_34_17_n_1310 = ~mul_34_17_n_1309;
 assign mul_34_17_n_1306 = ~mul_34_17_n_1305;
 assign mul_34_17_n_1294 = ~mul_34_17_n_1293;
 assign mul_34_17_n_1292 = ~mul_34_17_n_1291;
 assign mul_34_17_n_1286 = ~mul_34_17_n_1285;
 assign mul_34_17_n_1280 = ~mul_34_17_n_1279;
 assign mul_34_17_n_1270 = ~mul_34_17_n_1269;
 assign mul_34_17_n_1265 = ~mul_34_17_n_1264;
 assign mul_34_17_n_1260 = ~mul_34_17_n_1259;
 assign mul_34_17_n_1251 = ~mul_34_17_n_1250;
 assign mul_34_17_n_1244 = ~mul_34_17_n_1243;
 assign mul_34_17_n_1242 = ~mul_34_17_n_1241;
 assign mul_34_17_n_1237 = ~mul_34_17_n_1236;
 assign mul_34_17_n_1229 = ~mul_34_17_n_1228;
 assign mul_34_17_n_1223 = ~mul_34_17_n_1222;
 assign mul_34_17_n_1218 = ~mul_34_17_n_1217;
 assign mul_34_17_n_1216 = ~mul_34_17_n_1215;
 assign mul_34_17_n_1212 = ~mul_34_17_n_1211;
 assign mul_34_17_n_1210 = ~mul_34_17_n_1209;
 assign mul_34_17_n_1202 = ~mul_34_17_n_1201;
 assign mul_34_17_n_1199 = ~mul_34_17_n_1198;
 assign mul_34_17_n_1197 = ~mul_34_17_n_1196;
 assign mul_34_17_n_1195 = ~mul_34_17_n_1194;
 assign mul_34_17_n_1193 = ~mul_34_17_n_1192;
 assign mul_34_17_n_1191 = ~mul_34_17_n_1190;
 assign mul_34_17_n_1189 = ~mul_34_17_n_1188;
 assign mul_34_17_n_1184 = ~mul_34_17_n_1183;
 assign mul_34_17_n_1179 = ~mul_34_17_n_1178;
 assign mul_34_17_n_1176 = ~mul_34_17_n_1175;
 assign mul_34_17_n_1165 = ~mul_34_17_n_1164;
 assign mul_34_17_n_1163 = ~mul_34_17_n_1162;
 assign mul_34_17_n_1160 = ~mul_34_17_n_1159;
 assign mul_34_17_n_1157 = ~mul_34_17_n_1156;
 assign mul_34_17_n_1155 = ~mul_34_17_n_1154;
 assign mul_34_17_n_1146 = ~mul_34_17_n_1145;
 assign mul_34_17_n_1138 = ~mul_34_17_n_1137;
 assign mul_34_17_n_1136 = ~mul_34_17_n_1135;
 assign mul_34_17_n_1130 = ~mul_34_17_n_1129;
 assign mul_34_17_n_1127 = ~mul_34_17_n_1126;
 assign mul_34_17_n_1125 = ~mul_34_17_n_1124;
 assign mul_34_17_n_1123 = ~mul_34_17_n_1122;
 assign mul_34_17_n_1116 = ~mul_34_17_n_1115;
 assign mul_34_17_n_1113 = ~mul_34_17_n_1112;
 assign mul_34_17_n_1110 = ~mul_34_17_n_1109;
 assign mul_34_17_n_1104 = ~mul_34_17_n_1103;
 assign mul_34_17_n_1101 = ~mul_34_17_n_1100;
 assign mul_34_17_n_1098 = ~mul_34_17_n_1097;
 assign mul_34_17_n_1095 = ~mul_34_17_n_1094;
 assign mul_34_17_n_1093 = ~mul_34_17_n_1092;
 assign mul_34_17_n_1089 = ~mul_34_17_n_1088;
 assign mul_34_17_n_1085 = ~mul_34_17_n_1084;
 assign mul_34_17_n_1078 = ~mul_34_17_n_1077;
 assign mul_34_17_n_1075 = ~mul_34_17_n_1074;
 assign mul_34_17_n_1071 = ~mul_34_17_n_1070;
 assign mul_34_17_n_1065 = ~mul_34_17_n_1064;
 assign mul_34_17_n_1058 = ~mul_34_17_n_1057;
 assign mul_34_17_n_1046 = ~mul_34_17_n_1045;
 assign mul_34_17_n_1043 = ~mul_34_17_n_1042;
 assign mul_34_17_n_1038 = ~mul_34_17_n_1037;
 assign mul_34_17_n_1033 = ~mul_34_17_n_1032;
 assign mul_34_17_n_1031 = ~mul_34_17_n_1030;
 assign mul_34_17_n_1029 = ~mul_34_17_n_1028;
 assign mul_34_17_n_1025 = ~mul_34_17_n_1024;
 assign mul_34_17_n_1022 = ~mul_34_17_n_1021;
 assign mul_34_17_n_1016 = ~mul_34_17_n_1015;
 assign mul_34_17_n_1008 = ~mul_34_17_n_1007;
 assign mul_34_17_n_993 = ~mul_34_17_n_992;
 assign mul_34_17_n_980 = ~mul_34_17_n_979;
 assign mul_34_17_n_975 = ~mul_34_17_n_974;
 assign mul_34_17_n_972 = ~mul_34_17_n_971;
 assign mul_34_17_n_970 = ~mul_34_17_n_969;
 assign mul_34_17_n_966 = ~mul_34_17_n_965;
 assign mul_34_17_n_963 = ~mul_34_17_n_962;
 assign mul_34_17_n_960 = ~mul_34_17_n_959;
 assign mul_34_17_n_957 = ~mul_34_17_n_956;
 assign mul_34_17_n_954 = ~mul_34_17_n_953;
 assign mul_34_17_n_948 = ~mul_34_17_n_947;
 assign mul_34_17_n_942 = ~mul_34_17_n_941;
 assign mul_34_17_n_935 = ~mul_34_17_n_934;
 assign mul_34_17_n_930 = ~mul_34_17_n_929;
 assign mul_34_17_n_922 = ~mul_34_17_n_921;
 assign mul_34_17_n_919 = ~mul_34_17_n_918;
 assign mul_34_17_n_914 = ~mul_34_17_n_913;
 assign mul_34_17_n_907 = ~mul_34_17_n_906;
 assign mul_34_17_n_901 = ~mul_34_17_n_900;
 assign mul_34_17_n_898 = ~mul_34_17_n_897;
 assign mul_34_17_n_886 = ~mul_34_17_n_885;
 assign mul_34_17_n_883 = ~mul_34_17_n_882;
 assign mul_34_17_n_880 = ~mul_34_17_n_879;
 assign mul_34_17_n_875 = ~mul_34_17_n_874;
 assign mul_34_17_n_873 = ~mul_34_17_n_872;
 assign mul_34_17_n_869 = ~mul_34_17_n_868;
 assign mul_34_17_n_863 = ~mul_34_17_n_862;
 assign mul_34_17_n_860 = ~mul_34_17_n_859;
 assign mul_34_17_n_858 = ~mul_34_17_n_857;
 assign mul_34_17_n_848 = ~mul_34_17_n_847;
 assign mul_34_17_n_841 = ~mul_34_17_n_840;
 assign mul_34_17_n_828 = ~mul_34_17_n_827;
 assign mul_34_17_n_798 = ~mul_34_17_n_797;
 assign mul_34_17_n_787 = ~mul_34_17_n_786;
 assign mul_34_17_n_785 = ~mul_34_17_n_784;
 assign mul_34_17_n_783 = ~mul_34_17_n_782;
 assign mul_34_17_n_780 = ~mul_34_17_n_779;
 assign mul_34_17_n_776 = ~mul_34_17_n_775;
 assign mul_34_17_n_774 = ~mul_34_17_n_773;
 assign mul_34_17_n_771 = ~mul_34_17_n_770;
 assign mul_34_17_n_767 = ~mul_34_17_n_766;
 assign mul_34_17_n_764 = ~mul_34_17_n_763;
 assign mul_34_17_n_762 = ~mul_34_17_n_761;
 assign mul_34_17_n_760 = ~mul_34_17_n_759;
 assign mul_34_17_n_758 = ~mul_34_17_n_757;
 assign mul_34_17_n_756 = ~mul_34_17_n_755;
 assign mul_34_17_n_749 = ~mul_34_17_n_748;
 assign mul_34_17_n_746 = ~mul_34_17_n_745;
 assign mul_34_17_n_742 = ~mul_34_17_n_741;
 assign mul_34_17_n_737 = ~mul_34_17_n_736;
 assign mul_34_17_n_729 = ~mul_34_17_n_728;
 assign mul_34_17_n_720 = ~mul_34_17_n_719;
 assign mul_34_17_n_717 = ~mul_34_17_n_716;
 assign mul_34_17_n_690 = ~mul_34_17_n_691;
 assign mul_34_17_n_688 = ~mul_34_17_n_689;
 assign mul_34_17_n_686 = ~mul_34_17_n_687;
 assign mul_34_17_n_684 = ~mul_34_17_n_685;
 assign mul_34_17_n_682 = ~mul_34_17_n_683;
 assign mul_34_17_n_680 = ~mul_34_17_n_681;
 assign mul_34_17_n_678 = ~mul_34_17_n_679;
 assign mul_34_17_n_676 = ~mul_34_17_n_677;
 assign mul_34_17_n_674 = ~mul_34_17_n_675;
 assign mul_34_17_n_672 = ~mul_34_17_n_673;
 assign mul_34_17_n_670 = ~mul_34_17_n_671;
 assign mul_34_17_n_668 = ~mul_34_17_n_669;
 assign mul_34_17_n_666 = ~mul_34_17_n_667;
 assign mul_34_17_n_664 = ~mul_34_17_n_665;
 assign mul_34_17_n_662 = ~mul_34_17_n_663;
 assign mul_34_17_n_660 = ~mul_34_17_n_661;
 assign mul_34_17_n_658 = ~mul_34_17_n_659;
 assign mul_34_17_n_656 = ~mul_34_17_n_657;
 assign mul_34_17_n_654 = ~mul_34_17_n_655;
 assign mul_34_17_n_653 = ({in2[25]} ^ {in1[61]});
 assign mul_34_17_n_652 = ~({in2[61]} ^ {in1[25]});
 assign mul_34_17_n_651 = ~({in2[27]} ^ {in1[59]});
 assign mul_34_17_n_650 = ({in2[59]} ^ {in1[27]});
 assign mul_34_17_n_649 = ({in2[29]} ^ {in1[57]});
 assign mul_34_17_n_648 = ({in2[31]} ^ {in1[55]});
 assign mul_34_17_n_647 = ({in2[33]} ^ {in1[53]});
 assign mul_34_17_n_646 = ({in2[35]} ^ {in1[51]});
 assign mul_34_17_n_645 = ({in2[37]} ^ {in1[49]});
 assign mul_34_17_n_644 = ({in2[39]} ^ {in1[47]});
 assign mul_34_17_n_643 = ({in2[41]} ^ {in1[45]});
 assign mul_34_17_n_642 = ({in2[43]} ^ {in1[43]});
 assign mul_34_17_n_641 = ({in2[45]} ^ {in1[41]});
 assign mul_34_17_n_640 = ({in2[47]} ^ {in1[39]});
 assign mul_34_17_n_639 = ({in2[49]} ^ {in1[37]});
 assign mul_34_17_n_638 = ({in2[51]} ^ {in1[35]});
 assign mul_34_17_n_637 = ({in2[53]} ^ {in1[33]});
 assign mul_34_17_n_636 = ~({in2[55]} ^ {in1[31]});
 assign mul_34_17_n_635 = ({in2[57]} ^ {in1[29]});
 assign mul_34_17_n_634 = ({in2[63]} ^ {in1[23]});
 assign mul_34_17_n_1687 = ~({in2[25]} ^ {in1[21]});
 assign mul_34_17_n_1686 = ~({in2[25]} ^ {in1[46]});
 assign mul_34_17_n_1684 = ~({in2[25]} ^ {in1[56]});
 assign mul_34_17_n_1683 = ({in2[25]} ^ {in1[17]});
 assign mul_34_17_n_1681 = ~({in2[25]} ^ {in1[52]});
 assign mul_34_17_n_1680 = ({in2[25]} ^ {in1[60]});
 assign mul_34_17_n_1678 = ~({in2[25]} ^ {in1[43]});
 assign mul_34_17_n_1677 = ~({in2[25]} ^ {in1[20]});
 assign mul_34_17_n_1675 = ~({in2[25]} ^ {in1[47]});
 assign mul_34_17_n_1673 = ~({in2[25]} ^ {in1[3]});
 assign mul_34_17_n_1671 = ({in2[25]} ^ {in1[18]});
 assign mul_34_17_n_1670 = ~({in2[25]} ^ {in1[22]});
 assign mul_34_17_n_1669 = ~({in2[25]} ^ {in1[24]});
 assign mul_34_17_n_1667 = ~({in2[25]} ^ {in1[13]});
 assign mul_34_17_n_1665 = ~({in2[25]} ^ {in1[57]});
 assign mul_34_17_n_1664 = ({in2[27]} ^ {in1[55]});
 assign mul_34_17_n_1663 = ({in2[27]} ^ {in1[54]});
 assign mul_34_17_n_1662 = ({in2[27]} ^ {in1[28]});
 assign mul_34_17_n_1661 = ({in2[27]} ^ {in1[29]});
 assign mul_34_17_n_1660 = ({in2[27]} ^ {in1[51]});
 assign mul_34_17_n_1659 = ~({in2[27]} ^ {in1[5]});
 assign mul_34_17_n_1657 = ~({in2[27]} ^ {in1[26]});
 assign mul_34_17_n_1655 = ~({in2[27]} ^ {in1[13]});
 assign mul_34_17_n_1654 = ({in2[27]} ^ {in1[30]});
 assign mul_34_17_n_1652 = ~({in2[27]} ^ {in1[36]});
 assign mul_34_17_n_1651 = ~({in2[27]} ^ {in1[22]});
 assign mul_34_17_n_1649 = ~({in2[27]} ^ {in1[40]});
 assign mul_34_17_n_1648 = ({in2[27]} ^ {in1[41]});
 assign mul_34_17_n_1647 = ~({in2[27]} ^ {in1[43]});
 assign mul_34_17_n_1646 = ({in2[27]} ^ {in1[56]});
 assign mul_34_17_n_1645 = ~({in2[27]} ^ {in1[14]});
 assign mul_34_17_n_1644 = ~({in2[27]} ^ {in1[39]});
 assign mul_34_17_n_1643 = ~({in2[27]} ^ {in1[44]});
 assign mul_34_17_n_1642 = ({in2[27]} ^ {in1[49]});
 assign mul_34_17_n_1640 = ~({in2[27]} ^ {in1[37]});
 assign mul_34_17_n_1639 = ({in2[27]} ^ {in1[57]});
 assign mul_34_17_n_1638 = ~({in2[27]} ^ {in1[21]});
 assign mul_34_17_n_1636 = ~({in2[27]} ^ {in1[31]});
 assign mul_34_17_n_1634 = ({in2[27]} ^ {in1[48]});
 assign mul_34_17_n_1633 = ({in2[27]} ^ {in1[3]});
 assign mul_34_17_n_1632 = ({in2[25]} ^ {in1[42]});
 assign mul_34_17_n_1631 = ~({in2[27]} ^ {in1[24]});
 assign mul_34_17_n_1630 = ({in2[27]} ^ {in1[8]});
 assign mul_34_17_n_1629 = ~({in2[27]} ^ {in1[25]});
 assign mul_34_17_n_1628 = ({in2[27]} ^ {in1[10]});
 assign mul_34_17_n_1627 = ~({in2[27]} ^ {in1[15]});
 assign mul_34_17_n_1626 = ({in2[25]} ^ {in1[30]});
 assign mul_34_17_n_1624 = ({in2[27]} ^ {in1[6]});
 assign mul_34_17_n_1623 = ({in2[27]} ^ {in1[53]});
 assign mul_34_17_n_1622 = ({in2[27]} ^ {in1[52]});
 assign mul_34_17_n_1620 = ({in2[27]} ^ {in1[58]});
 assign mul_34_17_n_1619 = ({in2[27]} ^ {in1[34]});
 assign mul_34_17_n_1617 = ~({in2[27]} ^ {in1[4]});
 assign mul_34_17_n_1616 = ~({in2[27]} ^ {in1[47]});
 assign mul_34_17_n_1615 = ~({in2[27]} ^ {in1[19]});
 assign mul_34_17_n_1614 = ~({in2[27]} ^ {in1[46]});
 assign mul_34_17_n_1612 = ~({in2[27]} ^ {in1[33]});
 assign mul_34_17_n_1611 = ~({in2[27]} ^ {in1[18]});
 assign mul_34_17_n_1609 = ~({in2[27]} ^ {in1[2]});
 assign mul_34_17_n_1607 = ~({in2[27]} ^ {in1[1]});
 assign mul_34_17_n_1606 = ({in2[27]} ^ {in1[11]});
 assign mul_34_17_n_1605 = ({in2[27]} ^ {in1[12]});
 assign mul_34_17_n_1603 = ~({in2[27]} ^ {in1[35]});
 assign mul_34_17_n_1601 = ~({in2[27]} ^ {in1[42]});
 assign mul_34_17_n_1600 = ~({in2[27]} ^ {in1[17]});
 assign mul_34_17_n_1599 = ~({in2[27]} ^ {in1[32]});
 assign mul_34_17_n_1598 = ~({in2[27]} ^ {in1[16]});
 assign mul_34_17_n_1597 = ({in2[27]} ^ {in1[50]});
 assign mul_34_17_n_1596 = ~({in2[27]} ^ {in1[23]});
 assign mul_34_17_n_1595 = ({in2[27]} ^ {in1[27]});
 assign mul_34_17_n_1594 = ~({in2[27]} ^ {in1[45]});
 assign mul_34_17_n_1593 = ({in2[27]} ^ {in1[7]});
 assign mul_34_17_n_1592 = ({in2[27]} ^ {in1[9]});
 assign mul_34_17_n_1591 = ~({in2[27]} ^ {in1[20]});
 assign mul_34_17_n_1590 = ~({in2[27]} ^ {in1[38]});
 assign mul_34_17_n_1589 = ({in2[59]} ^ {in1[24]});
 assign mul_34_17_n_1587 = ~({in2[29]} ^ {in1[52]});
 assign mul_34_17_n_1586 = ({in2[29]} ^ {in1[54]});
 assign mul_34_17_n_1585 = ({in2[29]} ^ {in1[5]});
 assign mul_34_17_n_1584 = ({in2[29]} ^ {in1[36]});
 assign mul_34_17_n_1583 = ({in2[29]} ^ {in1[56]});
 assign mul_34_17_n_1581 = ~({in2[29]} ^ {in1[46]});
 assign mul_34_17_n_1579 = ~({in2[29]} ^ {in1[14]});
 assign mul_34_17_n_1578 = ({in2[29]} ^ {in1[55]});
 assign mul_34_17_n_1577 = ({in2[29]} ^ {in1[6]});
 assign mul_34_17_n_1576 = ~({in2[25]} ^ {in1[51]});
 assign mul_34_17_n_1575 = ~({in2[29]} ^ {in1[3]});
 assign mul_34_17_n_1574 = ({in2[29]} ^ {in1[8]});
 assign mul_34_17_n_1573 = ({in2[29]} ^ {in1[23]});
 assign mul_34_17_n_1572 = ({in2[29]} ^ {in1[31]});
 assign mul_34_17_n_1571 = ({in2[29]} ^ {in1[32]});
 assign mul_34_17_n_1570 = ~({in2[29]} ^ {in1[18]});
 assign mul_34_17_n_1569 = ({in2[29]} ^ {in1[33]});
 assign mul_34_17_n_1568 = ~({in2[29]} ^ {in1[49]});
 assign mul_34_17_n_1567 = ({in2[29]} ^ {in1[28]});
 assign mul_34_17_n_1566 = ~({in2[29]} ^ {in1[10]});
 assign mul_34_17_n_1565 = ~({in2[29]} ^ {in1[16]});
 assign mul_34_17_n_1563 = ~({in2[29]} ^ {in1[2]});
 assign mul_34_17_n_1562 = ~({in2[29]} ^ {in1[20]});
 assign mul_34_17_n_1561 = ({in2[29]} ^ {in1[38]});
 assign mul_34_17_n_1560 = ({in2[29]} ^ {in1[24]});
 assign mul_34_17_n_1559 = ({in2[29]} ^ {in1[29]});
 assign mul_34_17_n_1558 = ({in2[29]} ^ {in1[37]});
 assign mul_34_17_n_1556 = ({in2[29]} ^ {in1[9]});
 assign mul_34_17_n_1555 = ({in2[29]} ^ {in1[25]});
 assign mul_34_17_n_1553 = ~({in2[29]} ^ {in1[12]});
 assign mul_34_17_n_1551 = ~({in2[29]} ^ {in1[50]});
 assign mul_34_17_n_1550 = ({in2[29]} ^ {in1[26]});
 assign mul_34_17_n_1549 = ~({in2[29]} ^ {in1[11]});
 assign mul_34_17_n_1548 = ({in2[29]} ^ {in1[30]});
 assign mul_34_17_n_1546 = ~({in2[29]} ^ {in1[48]});
 assign mul_34_17_n_1545 = ~({in2[29]} ^ {in1[41]});
 assign mul_34_17_n_1544 = ~({in2[29]} ^ {in1[21]});
 assign mul_34_17_n_1543 = ({in2[29]} ^ {in1[51]});
 assign mul_34_17_n_1542 = ~({in2[29]} ^ {in1[19]});
 assign mul_34_17_n_1541 = ({in2[29]} ^ {in1[7]});
 assign mul_34_17_n_1539 = ~({in2[29]} ^ {in1[22]});
 assign mul_34_17_n_1537 = ~({in2[29]} ^ {in1[39]});
 assign mul_34_17_n_1536 = ~({in2[29]} ^ {in1[15]});
 assign mul_34_17_n_1535 = ({in2[29]} ^ {in1[13]});
 assign mul_34_17_n_1534 = ~({in2[29]} ^ {in1[42]});
 assign mul_34_17_n_1532 = ~({in2[29]} ^ {in1[53]});
 assign mul_34_17_n_1531 = ~({in2[29]} ^ {in1[17]});
 assign mul_34_17_n_1530 = ~({in2[29]} ^ {in1[40]});
 assign mul_34_17_n_1529 = ~({in2[29]} ^ {in1[44]});
 assign mul_34_17_n_1527 = ~({in2[29]} ^ {in1[4]});
 assign mul_34_17_n_1526 = ({in2[29]} ^ {in1[27]});
 assign mul_34_17_n_1525 = ({in2[29]} ^ {in1[47]});
 assign mul_34_17_n_1524 = ~({in2[29]} ^ {in1[43]});
 assign mul_34_17_n_1523 = ({in2[29]} ^ {in1[35]});
 assign mul_34_17_n_1522 = ~({in2[29]} ^ {in1[45]});
 assign mul_34_17_n_1521 = ({in2[29]} ^ {in1[1]});
 assign mul_34_17_n_1520 = ({in2[29]} ^ {in1[34]});
 assign mul_34_17_n_1519 = ~({in2[61]} ^ {in1[24]});
 assign mul_34_17_n_1517 = ~({in2[31]} ^ {in1[49]});
 assign mul_34_17_n_1515 = ~({in2[31]} ^ {in1[10]});
 assign mul_34_17_n_1514 = ({in2[31]} ^ {in1[54]});
 assign mul_34_17_n_1513 = ({in2[31]} ^ {in1[37]});
 assign mul_34_17_n_1512 = ({in2[31]} ^ {in1[1]});
 assign mul_34_17_n_1510 = ~({in2[31]} ^ {in1[28]});
 assign mul_34_17_n_1509 = ({in2[31]} ^ {in1[23]});
 assign mul_34_17_n_1507 = ({in2[31]} ^ {in1[5]});
 assign mul_34_17_n_1506 = ({in2[31]} ^ {in1[25]});
 assign mul_34_17_n_1505 = ~({in2[31]} ^ {in1[18]});
 assign mul_34_17_n_1503 = ~({in2[31]} ^ {in1[52]});
 assign mul_34_17_n_1501 = ~({in2[31]} ^ {in1[46]});
 assign mul_34_17_n_1500 = ~({in2[31]} ^ {in1[7]});
 assign mul_34_17_n_1498 = ~({in2[31]} ^ {in1[22]});
 assign mul_34_17_n_1497 = ({in2[31]} ^ {in1[20]});
 assign mul_34_17_n_1496 = ~({in2[31]} ^ {in1[17]});
 assign mul_34_17_n_1495 = ({in2[31]} ^ {in1[33]});
 assign mul_34_17_n_1493 = ~({in2[31]} ^ {in1[38]});
 assign mul_34_17_n_1491 = ~({in2[31]} ^ {in1[41]});
 assign mul_34_17_n_1489 = ~({in2[31]} ^ {in1[51]});
 assign mul_34_17_n_1488 = ~({in2[31]} ^ {in1[30]});
 assign mul_34_17_n_1486 = ~({in2[31]} ^ {in1[21]});
 assign mul_34_17_n_1485 = ~({in2[31]} ^ {in1[31]});
 assign mul_34_17_n_1483 = ~({in2[31]} ^ {in1[42]});
 assign mul_34_17_n_1482 = ({in2[31]} ^ {in1[3]});
 assign mul_34_17_n_1481 = ~({in2[31]} ^ {in1[16]});
 assign mul_34_17_n_1480 = ({in2[31]} ^ {in1[34]});
 assign mul_34_17_n_1479 = ({in2[31]} ^ {in1[4]});
 assign mul_34_17_n_1478 = ~({in2[31]} ^ {in1[45]});
 assign mul_34_17_n_1477 = ({in2[31]} ^ {in1[35]});
 assign mul_34_17_n_1476 = ~({in2[25]} ^ {in1[39]});
 assign mul_34_17_n_1474 = ~({in2[31]} ^ {in1[47]});
 assign mul_34_17_n_1473 = ~({in2[31]} ^ {in1[44]});
 assign mul_34_17_n_1472 = ({in2[31]} ^ {in1[11]});
 assign mul_34_17_n_1471 = ~({in2[31]} ^ {in1[40]});
 assign mul_34_17_n_1469 = ~({in2[31]} ^ {in1[12]});
 assign mul_34_17_n_1468 = ~({in2[31]} ^ {in1[43]});
 assign mul_34_17_n_1467 = ~({in2[31]} ^ {in1[8]});
 assign mul_34_17_n_1466 = ~({in2[31]} ^ {in1[29]});
 assign mul_34_17_n_1464 = ({in2[31]} ^ {in1[19]});
 assign mul_34_17_n_1463 = ~({in2[31]} ^ {in1[9]});
 assign mul_34_17_n_1461 = ~({in2[31]} ^ {in1[15]});
 assign mul_34_17_n_1460 = ({in2[31]} ^ {in1[36]});
 assign mul_34_17_n_1459 = ({in2[31]} ^ {in1[53]});
 assign mul_34_17_n_1458 = ({in2[31]} ^ {in1[27]});
 assign mul_34_17_n_1457 = ~({in2[31]} ^ {in1[48]});
 assign mul_34_17_n_1456 = ({in2[31]} ^ {in1[2]});
 assign mul_34_17_n_1454 = ~({in2[31]} ^ {in1[32]});
 assign mul_34_17_n_1453 = ({in2[31]} ^ {in1[50]});
 assign mul_34_17_n_1452 = ({in2[31]} ^ {in1[26]});
 assign mul_34_17_n_1451 = ~({in2[31]} ^ {in1[39]});
 assign mul_34_17_n_1450 = ~({in2[31]} ^ {in1[6]});
 assign mul_34_17_n_1449 = ~({in2[31]} ^ {in1[13]});
 assign mul_34_17_n_1448 = ({in2[31]} ^ {in1[24]});
 assign mul_34_17_n_1446 = ~({in2[31]} ^ {in1[14]});
 assign mul_34_17_n_1444 = ~({in2[33]} ^ {in1[47]});
 assign mul_34_17_n_1443 = ~({in2[33]} ^ {in1[39]});
 assign mul_34_17_n_1442 = ({in2[33]} ^ {in1[21]});
 assign mul_34_17_n_1441 = ({in2[33]} ^ {in1[50]});
 assign mul_34_17_n_1439 = ({in2[33]} ^ {in1[10]});
 assign mul_34_17_n_1438 = ({in2[33]} ^ {in1[16]});
 assign mul_34_17_n_1437 = ({in2[33]} ^ {in1[51]});
 assign mul_34_17_n_1436 = ({in2[33]} ^ {in1[52]});
 assign mul_34_17_n_1435 = ({in2[33]} ^ {in1[18]});
 assign mul_34_17_n_1434 = ({in2[33]} ^ {in1[35]});
 assign mul_34_17_n_1432 = ~({in2[33]} ^ {in1[46]});
 assign mul_34_17_n_1430 = ~({in2[33]} ^ {in1[32]});
 assign mul_34_17_n_1429 = ({in2[33]} ^ {in1[6]});
 assign mul_34_17_n_1428 = ({in2[33]} ^ {in1[2]});
 assign mul_34_17_n_1427 = ({in2[33]} ^ {in1[25]});
 assign mul_34_17_n_1426 = ({in2[33]} ^ {in1[44]});
 assign mul_34_17_n_1424 = ~({in2[33]} ^ {in1[3]});
 assign mul_34_17_n_1423 = ({in2[33]} ^ {in1[13]});
 assign mul_34_17_n_1422 = ({in2[33]} ^ {in1[43]});
 assign mul_34_17_n_1420 = ~({in2[33]} ^ {in1[14]});
 assign mul_34_17_n_1419 = ({in2[33]} ^ {in1[34]});
 assign mul_34_17_n_1417 = ~({in2[33]} ^ {in1[15]});
 assign mul_34_17_n_1415 = ({in2[33]} ^ {in1[12]});
 assign mul_34_17_n_1414 = ({in2[25]} ^ {in1[8]});
 assign mul_34_17_n_1413 = ({in2[33]} ^ {in1[20]});
 assign mul_34_17_n_1412 = ~({in2[33]} ^ {in1[27]});
 assign mul_34_17_n_1411 = ~({in2[33]} ^ {in1[28]});
 assign mul_34_17_n_1410 = ({in2[33]} ^ {in1[22]});
 assign mul_34_17_n_1409 = ({in2[33]} ^ {in1[19]});
 assign mul_34_17_n_1407 = ~({in2[33]} ^ {in1[30]});
 assign mul_34_17_n_1405 = ~({in2[33]} ^ {in1[48]});
 assign mul_34_17_n_1403 = ~({in2[33]} ^ {in1[49]});
 assign mul_34_17_n_1401 = ~({in2[33]} ^ {in1[42]});
 assign mul_34_17_n_1399 = ~({in2[33]} ^ {in1[8]});
 assign mul_34_17_n_1398 = ~({in2[33]} ^ {in1[11]});
 assign mul_34_17_n_1397 = ({in2[33]} ^ {in1[33]});
 assign mul_34_17_n_1396 = ({in2[33]} ^ {in1[9]});
 assign mul_34_17_n_1395 = ~({in2[33]} ^ {in1[37]});
 assign mul_34_17_n_1393 = ~({in2[33]} ^ {in1[31]});
 assign mul_34_17_n_1392 = ~({in2[33]} ^ {in1[29]});
 assign mul_34_17_n_1391 = ({in2[33]} ^ {in1[23]});
 assign mul_34_17_n_1390 = ({in2[33]} ^ {in1[24]});
 assign mul_34_17_n_1389 = ~({in2[33]} ^ {in1[38]});
 assign mul_34_17_n_1387 = ~({in2[33]} ^ {in1[5]});
 assign mul_34_17_n_1386 = ({in2[33]} ^ {in1[17]});
 assign mul_34_17_n_1385 = ({in2[59]} ^ {in1[25]});
 assign mul_34_17_n_1384 = ({in2[33]} ^ {in1[45]});
 assign mul_34_17_n_1382 = ~({in2[33]} ^ {in1[26]});
 assign mul_34_17_n_1381 = ~({in2[33]} ^ {in1[41]});
 assign mul_34_17_n_1379 = ~({in2[33]} ^ {in1[7]});
 assign mul_34_17_n_1378 = ~({in2[33]} ^ {in1[40]});
 assign mul_34_17_n_1376 = ~({in2[33]} ^ {in1[36]});
 assign mul_34_17_n_1375 = ~({in2[33]} ^ {in1[4]});
 assign mul_34_17_n_1374 = ({in2[33]} ^ {in1[1]});
 assign mul_34_17_n_1373 = ~({in2[35]} ^ {in1[3]});
 assign mul_34_17_n_1372 = ({in2[35]} ^ {in1[1]});
 assign mul_34_17_n_1370 = ~({in2[35]} ^ {in1[28]});
 assign mul_34_17_n_1369 = ({in2[35]} ^ {in1[22]});
 assign mul_34_17_n_1368 = ~({in2[35]} ^ {in1[13]});
 assign mul_34_17_n_1367 = ({in2[35]} ^ {in1[21]});
 assign mul_34_17_n_1366 = ({in2[35]} ^ {in1[30]});
 assign mul_34_17_n_1364 = ({in2[35]} ^ {in1[38]});
 assign mul_34_17_n_1363 = ~({in2[35]} ^ {in1[12]});
 assign mul_34_17_n_1362 = ({in2[35]} ^ {in1[45]});
 assign mul_34_17_n_1360 = ({in2[35]} ^ {in1[2]});
 assign mul_34_17_n_1358 = ~({in2[35]} ^ {in1[9]});
 assign mul_34_17_n_1357 = ({in2[35]} ^ {in1[29]});
 assign mul_34_17_n_1356 = ~({in2[35]} ^ {in1[39]});
 assign mul_34_17_n_1355 = ~({in2[35]} ^ {in1[14]});
 assign mul_34_17_n_1354 = ({in2[35]} ^ {in1[32]});
 assign mul_34_17_n_1353 = ~({in2[35]} ^ {in1[40]});
 assign mul_34_17_n_1352 = ({in2[35]} ^ {in1[17]});
 assign mul_34_17_n_1351 = ({in2[35]} ^ {in1[19]});
 assign mul_34_17_n_1350 = ({in2[35]} ^ {in1[48]});
 assign mul_34_17_n_1349 = ~({in2[35]} ^ {in1[27]});
 assign mul_34_17_n_1348 = ~({in2[35]} ^ {in1[8]});
 assign mul_34_17_n_1347 = ~({in2[35]} ^ {in1[35]});
 assign mul_34_17_n_1345 = ~({in2[35]} ^ {in1[10]});
 assign mul_34_17_n_1344 = ({in2[35]} ^ {in1[37]});
 assign mul_34_17_n_1343 = ({in2[35]} ^ {in1[20]});
 assign mul_34_17_n_1342 = ~({in2[25]} ^ {in1[40]});
 assign mul_34_17_n_1341 = ~({in2[35]} ^ {in1[34]});
 assign mul_34_17_n_1340 = ({in2[35]} ^ {in1[16]});
 assign mul_34_17_n_1338 = ({in2[35]} ^ {in1[41]});
 assign mul_34_17_n_1337 = ({in2[59]} ^ {in1[26]});
 assign mul_34_17_n_1335 = ~({in2[35]} ^ {in1[46]});
 assign mul_34_17_n_1333 = ~({in2[35]} ^ {in1[36]});
 assign mul_34_17_n_1332 = ({in2[35]} ^ {in1[31]});
 assign mul_34_17_n_1331 = ({in2[35]} ^ {in1[49]});
 assign mul_34_17_n_1330 = ({in2[35]} ^ {in1[43]});
 assign mul_34_17_n_1329 = ({in2[35]} ^ {in1[5]});
 assign mul_34_17_n_1328 = ({in2[35]} ^ {in1[50]});
 assign mul_34_17_n_1327 = ~({in2[35]} ^ {in1[26]});
 assign mul_34_17_n_1326 = ~({in2[35]} ^ {in1[25]});
 assign mul_34_17_n_1325 = ({in2[35]} ^ {in1[18]});
 assign mul_34_17_n_1323 = ~({in2[35]} ^ {in1[6]});
 assign mul_34_17_n_1322 = ({in2[35]} ^ {in1[42]});
 assign mul_34_17_n_1321 = ~({in2[35]} ^ {in1[11]});
 assign mul_34_17_n_1319 = ~({in2[35]} ^ {in1[47]});
 assign mul_34_17_n_1317 = ~({in2[35]} ^ {in1[15]});
 assign mul_34_17_n_1316 = ~({in2[35]} ^ {in1[7]});
 assign mul_34_17_n_1314 = ~({in2[35]} ^ {in1[33]});
 assign mul_34_17_n_1312 = ({in2[35]} ^ {in1[4]});
 assign mul_34_17_n_1311 = ({in2[35]} ^ {in1[23]});
 assign mul_34_17_n_1309 = ~({in2[35]} ^ {in1[24]});
 assign mul_34_17_n_1308 = ({in2[35]} ^ {in1[44]});
 assign mul_34_17_n_1307 = ~({in2[37]} ^ {in1[45]});
 assign mul_34_17_n_1305 = ~({in2[37]} ^ {in1[46]});
 assign mul_34_17_n_1304 = ~({in2[37]} ^ {in1[23]});
 assign mul_34_17_n_1303 = ~({in2[37]} ^ {in1[7]});
 assign mul_34_17_n_1302 = ~({in2[37]} ^ {in1[4]});
 assign mul_34_17_n_1301 = ({in2[37]} ^ {in1[30]});
 assign mul_34_17_n_1300 = ~({in2[37]} ^ {in1[6]});
 assign mul_34_17_n_1299 = ({in2[37]} ^ {in1[42]});
 assign mul_34_17_n_1298 = ({in2[37]} ^ {in1[17]});
 assign mul_34_17_n_1297 = ({in2[37]} ^ {in1[40]});
 assign mul_34_17_n_1296 = ~({in2[37]} ^ {in1[34]});
 assign mul_34_17_n_1295 = ~({in2[37]} ^ {in1[27]});
 assign mul_34_17_n_1293 = ~({in2[37]} ^ {in1[2]});
 assign mul_34_17_n_1291 = ~({in2[37]} ^ {in1[22]});
 assign mul_34_17_n_1290 = ({in2[37]} ^ {in1[21]});
 assign mul_34_17_n_1289 = ({in2[37]} ^ {in1[19]});
 assign mul_34_17_n_1288 = ~({in2[37]} ^ {in1[36]});
 assign mul_34_17_n_1287 = ({in2[37]} ^ {in1[14]});
 assign mul_34_17_n_1285 = ~({in2[37]} ^ {in1[44]});
 assign mul_34_17_n_1284 = ~({in2[37]} ^ {in1[35]});
 assign mul_34_17_n_1283 = ({in2[37]} ^ {in1[41]});
 assign mul_34_17_n_1282 = ~({in2[37]} ^ {in1[28]});
 assign mul_34_17_n_1281 = ~({in2[37]} ^ {in1[33]});
 assign mul_34_17_n_1279 = ~({in2[25]} ^ {in1[15]});
 assign mul_34_17_n_1278 = ~({in2[37]} ^ {in1[37]});
 assign mul_34_17_n_1277 = ({in2[37]} ^ {in1[20]});
 assign mul_34_17_n_1276 = ~({in2[37]} ^ {in1[26]});
 assign mul_34_17_n_1275 = ~({in2[37]} ^ {in1[10]});
 assign mul_34_17_n_1274 = ~({in2[37]} ^ {in1[3]});
 assign mul_34_17_n_1273 = ~({in2[37]} ^ {in1[8]});
 assign mul_34_17_n_1272 = ({in2[37]} ^ {in1[48]});
 assign mul_34_17_n_1271 = ~({in2[37]} ^ {in1[38]});
 assign mul_34_17_n_1269 = ({in2[37]} ^ {in1[29]});
 assign mul_34_17_n_1268 = ({in2[37]} ^ {in1[43]});
 assign mul_34_17_n_1267 = ~({in2[37]} ^ {in1[12]});
 assign mul_34_17_n_1266 = ~({in2[61]} ^ {in1[22]});
 assign mul_34_17_n_1264 = ~({in2[37]} ^ {in1[39]});
 assign mul_34_17_n_1263 = ({in2[37]} ^ {in1[1]});
 assign mul_34_17_n_1262 = ~({in2[37]} ^ {in1[5]});
 assign mul_34_17_n_1261 = ({in2[37]} ^ {in1[15]});
 assign mul_34_17_n_1259 = ({in2[37]} ^ {in1[13]});
 assign mul_34_17_n_1258 = ({in2[37]} ^ {in1[31]});
 assign mul_34_17_n_1257 = ({in2[37]} ^ {in1[47]});
 assign mul_34_17_n_1256 = ~({in2[37]} ^ {in1[25]});
 assign mul_34_17_n_1255 = ~({in2[37]} ^ {in1[9]});
 assign mul_34_17_n_1254 = ~({in2[37]} ^ {in1[24]});
 assign mul_34_17_n_1253 = ({in2[37]} ^ {in1[18]});
 assign mul_34_17_n_1252 = ~({in2[37]} ^ {in1[11]});
 assign mul_34_17_n_1250 = ~({in2[37]} ^ {in1[32]});
 assign mul_34_17_n_1249 = ({in2[37]} ^ {in1[16]});
 assign mul_34_17_n_1248 = ({in2[39]} ^ {in1[46]});
 assign mul_34_17_n_1247 = ({in2[39]} ^ {in1[25]});
 assign mul_34_17_n_1246 = ({in2[39]} ^ {in1[12]});
 assign mul_34_17_n_1245 = ({in2[39]} ^ {in1[13]});
 assign mul_34_17_n_1243 = ~({in2[39]} ^ {in1[40]});
 assign mul_34_17_n_1241 = ~({in2[39]} ^ {in1[15]});
 assign mul_34_17_n_1240 = ({in2[39]} ^ {in1[14]});
 assign mul_34_17_n_1239 = ~({in2[39]} ^ {in1[31]});
 assign mul_34_17_n_1238 = ~({in2[39]} ^ {in1[7]});
 assign mul_34_17_n_1236 = ~({in2[39]} ^ {in1[38]});
 assign mul_34_17_n_1235 = ~({in2[39]} ^ {in1[9]});
 assign mul_34_17_n_1234 = ~({in2[39]} ^ {in1[33]});
 assign mul_34_17_n_1233 = ({in2[25]} ^ {in1[5]});
 assign mul_34_17_n_1232 = ~({in2[39]} ^ {in1[10]});
 assign mul_34_17_n_1231 = ~({in2[39]} ^ {in1[37]});
 assign mul_34_17_n_1230 = ~({in2[39]} ^ {in1[30]});
 assign mul_34_17_n_1228 = ({in2[39]} ^ {in1[11]});
 assign mul_34_17_n_1227 = ~({in2[39]} ^ {in1[22]});
 assign mul_34_17_n_1226 = ~({in2[39]} ^ {in1[6]});
 assign mul_34_17_n_1225 = ~({in2[39]} ^ {in1[3]});
 assign mul_34_17_n_1224 = ({in2[39]} ^ {in1[44]});
 assign mul_34_17_n_1222 = ~({in2[39]} ^ {in1[1]});
 assign mul_34_17_n_1221 = ~({in2[39]} ^ {in1[36]});
 assign mul_34_17_n_1220 = ~({in2[39]} ^ {in1[2]});
 assign mul_34_17_n_1219 = ~({in2[39]} ^ {in1[16]});
 assign mul_34_17_n_1217 = ~({in2[39]} ^ {in1[17]});
 assign mul_34_17_n_1215 = ~({in2[39]} ^ {in1[5]});
 assign mul_34_17_n_1214 = ({in2[39]} ^ {in1[19]});
 assign mul_34_17_n_1213 = ~({in2[39]} ^ {in1[34]});
 assign mul_34_17_n_1211 = ~({in2[39]} ^ {in1[42]});
 assign mul_34_17_n_1209 = ~({in2[39]} ^ {in1[43]});
 assign mul_34_17_n_1208 = ~({in2[39]} ^ {in1[21]});
 assign mul_34_17_n_1207 = ~({in2[39]} ^ {in1[35]});
 assign mul_34_17_n_1206 = ({in2[39]} ^ {in1[39]});
 assign mul_34_17_n_1205 = ~({in2[39]} ^ {in1[23]});
 assign mul_34_17_n_1204 = ({in2[39]} ^ {in1[45]});
 assign mul_34_17_n_1203 = ~({in2[39]} ^ {in1[32]});
 assign mul_34_17_n_1201 = ~({in2[39]} ^ {in1[20]});
 assign mul_34_17_n_1200 = ~({in2[61]} ^ {in1[20]});
 assign mul_34_17_n_1198 = ~({in2[39]} ^ {in1[26]});
 assign mul_34_17_n_1196 = ~({in2[39]} ^ {in1[29]});
 assign mul_34_17_n_1194 = ~({in2[39]} ^ {in1[41]});
 assign mul_34_17_n_1192 = ~({in2[39]} ^ {in1[27]});
 assign mul_34_17_n_1190 = ({in2[39]} ^ {in1[4]});
 assign mul_34_17_n_1188 = ~({in2[39]} ^ {in1[24]});
 assign mul_34_17_n_1187 = ({in2[39]} ^ {in1[18]});
 assign mul_34_17_n_1186 = ({in2[39]} ^ {in1[28]});
 assign mul_34_17_n_1185 = ~({in2[39]} ^ {in1[8]});
 assign mul_34_17_n_1183 = ~({in2[41]} ^ {in1[2]});
 assign mul_34_17_n_1182 = ~({in2[41]} ^ {in1[10]});
 assign mul_34_17_n_1181 = ~({in2[41]} ^ {in1[14]});
 assign mul_34_17_n_1180 = ({in2[41]} ^ {in1[44]});
 assign mul_34_17_n_1178 = ~({in2[41]} ^ {in1[19]});
 assign mul_34_17_n_1177 = ({in2[41]} ^ {in1[16]});
 assign mul_34_17_n_1175 = ({in2[25]} ^ {in1[49]});
 assign mul_34_17_n_1174 = ~({in2[41]} ^ {in1[29]});
 assign mul_34_17_n_1173 = ~({in2[41]} ^ {in1[28]});
 assign mul_34_17_n_1172 = ~({in2[41]} ^ {in1[33]});
 assign mul_34_17_n_1171 = ~({in2[41]} ^ {in1[30]});
 assign mul_34_17_n_1170 = ~({in2[41]} ^ {in1[32]});
 assign mul_34_17_n_1169 = ({in2[41]} ^ {in1[39]});
 assign mul_34_17_n_1168 = ~({in2[41]} ^ {in1[6]});
 assign mul_34_17_n_1167 = ({in2[63]} ^ {in1[10]});
 assign mul_34_17_n_1166 = ({in2[41]} ^ {in1[24]});
 assign mul_34_17_n_1164 = ~({in2[41]} ^ {in1[5]});
 assign mul_34_17_n_1162 = ~({in2[41]} ^ {in1[17]});
 assign mul_34_17_n_1161 = ({in2[41]} ^ {in1[25]});
 assign mul_34_17_n_1159 = ~({in2[41]} ^ {in1[4]});
 assign mul_34_17_n_1158 = ({in2[41]} ^ {in1[23]});
 assign mul_34_17_n_1156 = ~({in2[41]} ^ {in1[26]});
 assign mul_34_17_n_1154 = ~({in2[41]} ^ {in1[12]});
 assign mul_34_17_n_1153 = ({in2[41]} ^ {in1[42]});
 assign mul_34_17_n_1152 = ({in2[41]} ^ {in1[40]});
 assign mul_34_17_n_1151 = ({in2[41]} ^ {in1[41]});
 assign mul_34_17_n_1150 = ~({in2[41]} ^ {in1[7]});
 assign mul_34_17_n_1149 = ~({in2[41]} ^ {in1[18]});
 assign mul_34_17_n_1148 = ({in2[41]} ^ {in1[38]});
 assign mul_34_17_n_1147 = ({in2[41]} ^ {in1[37]});
 assign mul_34_17_n_1145 = ({in2[41]} ^ {in1[35]});
 assign mul_34_17_n_1144 = ({in2[41]} ^ {in1[43]});
 assign mul_34_17_n_1143 = ~({in2[41]} ^ {in1[8]});
 assign mul_34_17_n_1142 = ~({in2[41]} ^ {in1[31]});
 assign mul_34_17_n_1141 = ({in2[41]} ^ {in1[20]});
 assign mul_34_17_n_1140 = ~({in2[41]} ^ {in1[11]});
 assign mul_34_17_n_1139 = ({in2[41]} ^ {in1[1]});
 assign mul_34_17_n_1137 = ~({in2[41]} ^ {in1[13]});
 assign mul_34_17_n_1135 = ~({in2[41]} ^ {in1[22]});
 assign mul_34_17_n_1134 = ~({in2[41]} ^ {in1[27]});
 assign mul_34_17_n_1133 = ~({in2[41]} ^ {in1[9]});
 assign mul_34_17_n_1132 = ({in2[41]} ^ {in1[36]});
 assign mul_34_17_n_1131 = ~({in2[41]} ^ {in1[3]});
 assign mul_34_17_n_1129 = ~({in2[41]} ^ {in1[21]});
 assign mul_34_17_n_1128 = ~({in2[41]} ^ {in1[34]});
 assign mul_34_17_n_1126 = ({in2[41]} ^ {in1[15]});
 assign mul_34_17_n_1124 = ~({in2[43]} ^ {in1[39]});
 assign mul_34_17_n_1122 = ({in2[43]} ^ {in1[18]});
 assign mul_34_17_n_1121 = ({in2[43]} ^ {in1[12]});
 assign mul_34_17_n_1120 = ({in2[43]} ^ {in1[41]});
 assign mul_34_17_n_1119 = ({in2[43]} ^ {in1[23]});
 assign mul_34_17_n_1118 = ({in2[43]} ^ {in1[13]});
 assign mul_34_17_n_1117 = ({in2[43]} ^ {in1[9]});
 assign mul_34_17_n_1115 = ~({in2[43]} ^ {in1[28]});
 assign mul_34_17_n_1114 = ({in2[43]} ^ {in1[37]});
 assign mul_34_17_n_1112 = ~({in2[59]} ^ {in1[18]});
 assign mul_34_17_n_1111 = ({in2[25]} ^ {in1[7]});
 assign mul_34_17_n_1109 = ~({in2[43]} ^ {in1[8]});
 assign mul_34_17_n_1108 = ({in2[43]} ^ {in1[11]});
 assign mul_34_17_n_1107 = ({in2[43]} ^ {in1[36]});
 assign mul_34_17_n_1106 = ({in2[43]} ^ {in1[6]});
 assign mul_34_17_n_1105 = ({in2[43]} ^ {in1[1]});
 assign mul_34_17_n_1103 = ~({in2[43]} ^ {in1[3]});
 assign mul_34_17_n_1102 = ({in2[43]} ^ {in1[10]});
 assign mul_34_17_n_1100 = ~({in2[43]} ^ {in1[20]});
 assign mul_34_17_n_1099 = ({in2[43]} ^ {in1[14]});
 assign mul_34_17_n_1097 = ~({in2[43]} ^ {in1[31]});
 assign mul_34_17_n_1096 = ({in2[43]} ^ {in1[42]});
 assign mul_34_17_n_1094 = ~({in2[43]} ^ {in1[38]});
 assign mul_34_17_n_1092 = ~({in2[43]} ^ {in1[26]});
 assign mul_34_17_n_1091 = ({in2[43]} ^ {in1[24]});
 assign mul_34_17_n_1090 = ~({in2[43]} ^ {in1[17]});
 assign mul_34_17_n_1088 = ~({in2[43]} ^ {in1[34]});
 assign mul_34_17_n_1087 = ({in2[43]} ^ {in1[30]});
 assign mul_34_17_n_1086 = ({in2[43]} ^ {in1[29]});
 assign mul_34_17_n_1084 = ~({in2[43]} ^ {in1[19]});
 assign mul_34_17_n_1083 = ({in2[43]} ^ {in1[5]});
 assign mul_34_17_n_1082 = ({in2[43]} ^ {in1[25]});
 assign mul_34_17_n_1081 = ~({in2[43]} ^ {in1[32]});
 assign mul_34_17_n_1080 = ({in2[43]} ^ {in1[35]});
 assign mul_34_17_n_1079 = ({in2[43]} ^ {in1[15]});
 assign mul_34_17_n_1077 = ~({in2[43]} ^ {in1[16]});
 assign mul_34_17_n_1076 = ({in2[43]} ^ {in1[22]});
 assign mul_34_17_n_1074 = ~({in2[43]} ^ {in1[4]});
 assign mul_34_17_n_1073 = ({in2[43]} ^ {in1[40]});
 assign mul_34_17_n_1072 = ({in2[43]} ^ {in1[21]});
 assign mul_34_17_n_1070 = ({in2[43]} ^ {in1[7]});
 assign mul_34_17_n_1069 = ~({in2[43]} ^ {in1[27]});
 assign mul_34_17_n_1068 = ~({in2[43]} ^ {in1[33]});
 assign mul_34_17_n_1067 = ({in2[43]} ^ {in1[2]});
 assign mul_34_17_n_1066 = ~({in2[45]} ^ {in1[37]});
 assign mul_34_17_n_1064 = ~({in2[45]} ^ {in1[36]});
 assign mul_34_17_n_1063 = ({in2[25]} ^ {in1[6]});
 assign mul_34_17_n_1062 = ({in2[45]} ^ {in1[21]});
 assign mul_34_17_n_1061 = ({in2[45]} ^ {in1[35]});
 assign mul_34_17_n_1060 = ({in2[45]} ^ {in1[10]});
 assign mul_34_17_n_1059 = ~({in2[45]} ^ {in1[29]});
 assign mul_34_17_n_1057 = ~({in2[63]} ^ {in1[6]});
 assign mul_34_17_n_1056 = ~({in2[45]} ^ {in1[26]});
 assign mul_34_17_n_1055 = ({in2[45]} ^ {in1[34]});
 assign mul_34_17_n_1054 = ({in2[45]} ^ {in1[11]});
 assign mul_34_17_n_1053 = ({in2[45]} ^ {in1[33]});
 assign mul_34_17_n_1052 = ~({in2[45]} ^ {in1[4]});
 assign mul_34_17_n_1051 = ({in2[45]} ^ {in1[39]});
 assign mul_34_17_n_1050 = ~({in2[45]} ^ {in1[31]});
 assign mul_34_17_n_1049 = ({in2[45]} ^ {in1[7]});
 assign mul_34_17_n_1048 = ~({in2[45]} ^ {in1[2]});
 assign mul_34_17_n_1047 = ({in2[45]} ^ {in1[22]});
 assign mul_34_17_n_1045 = ~({in2[45]} ^ {in1[17]});
 assign mul_34_17_n_1044 = ({in2[45]} ^ {in1[20]});
 assign mul_34_17_n_1042 = ~({in2[45]} ^ {in1[18]});
 assign mul_34_17_n_1041 = ~({in2[45]} ^ {in1[28]});
 assign mul_34_17_n_1040 = ({in2[45]} ^ {in1[12]});
 assign mul_34_17_n_1039 = ({in2[45]} ^ {in1[6]});
 assign mul_34_17_n_1037 = ~({in2[45]} ^ {in1[14]});
 assign mul_34_17_n_1036 = ({in2[45]} ^ {in1[23]});
 assign mul_34_17_n_1035 = ~({in2[45]} ^ {in1[15]});
 assign mul_34_17_n_1034 = ({in2[45]} ^ {in1[40]});
 assign mul_34_17_n_1032 = ~({in2[45]} ^ {in1[16]});
 assign mul_34_17_n_1030 = ~({in2[45]} ^ {in1[32]});
 assign mul_34_17_n_1028 = ~({in2[45]} ^ {in1[1]});
 assign mul_34_17_n_1027 = ~({in2[45]} ^ {in1[25]});
 assign mul_34_17_n_1026 = ~({in2[45]} ^ {in1[30]});
 assign mul_34_17_n_1024 = ~({in2[45]} ^ {in1[24]});
 assign mul_34_17_n_1023 = ~({in2[45]} ^ {in1[27]});
 assign mul_34_17_n_1021 = ~({in2[45]} ^ {in1[5]});
 assign mul_34_17_n_1020 = ({in2[45]} ^ {in1[9]});
 assign mul_34_17_n_1019 = ({in2[45]} ^ {in1[13]});
 assign mul_34_17_n_1018 = ({in2[45]} ^ {in1[19]});
 assign mul_34_17_n_1017 = ~({in2[45]} ^ {in1[3]});
 assign mul_34_17_n_1015 = ~({in2[45]} ^ {in1[38]});
 assign mul_34_17_n_1014 = ({in2[45]} ^ {in1[8]});
 assign mul_34_17_n_1013 = ~({in2[47]} ^ {in1[24]});
 assign mul_34_17_n_1012 = ({in2[47]} ^ {in1[5]});
 assign mul_34_17_n_1011 = ({in2[47]} ^ {in1[7]});
 assign mul_34_17_n_1010 = ({in2[47]} ^ {in1[38]});
 assign mul_34_17_n_1009 = ({in2[63]} ^ {in1[16]});
 assign mul_34_17_n_1007 = ~({in2[47]} ^ {in1[19]});
 assign mul_34_17_n_1006 = ~({in2[47]} ^ {in1[15]});
 assign mul_34_17_n_1005 = ~({in2[47]} ^ {in1[14]});
 assign mul_34_17_n_1004 = ~({in2[47]} ^ {in1[25]});
 assign mul_34_17_n_1003 = ({in2[25]} ^ {in1[27]});
 assign mul_34_17_n_1002 = ({in2[47]} ^ {in1[36]});
 assign mul_34_17_n_1001 = ({in2[47]} ^ {in1[28]});
 assign mul_34_17_n_1000 = ({in2[47]} ^ {in1[32]});
 assign mul_34_17_n_999 = ~({in2[47]} ^ {in1[16]});
 assign mul_34_17_n_998 = ({in2[47]} ^ {in1[31]});
 assign mul_34_17_n_997 = ({in2[47]} ^ {in1[11]});
 assign mul_34_17_n_996 = ({in2[47]} ^ {in1[33]});
 assign mul_34_17_n_995 = ({in2[47]} ^ {in1[10]});
 assign mul_34_17_n_994 = ({in2[47]} ^ {in1[37]});
 assign mul_34_17_n_992 = ~({in2[47]} ^ {in1[12]});
 assign mul_34_17_n_991 = ({in2[47]} ^ {in1[30]});
 assign mul_34_17_n_990 = ({in2[47]} ^ {in1[34]});
 assign mul_34_17_n_989 = ({in2[47]} ^ {in1[21]});
 assign mul_34_17_n_988 = ({in2[47]} ^ {in1[8]});
 assign mul_34_17_n_987 = ~({in2[47]} ^ {in1[17]});
 assign mul_34_17_n_986 = ({in2[47]} ^ {in1[1]});
 assign mul_34_17_n_985 = ~({in2[47]} ^ {in1[13]});
 assign mul_34_17_n_984 = ~({in2[47]} ^ {in1[23]});
 assign mul_34_17_n_983 = ({in2[47]} ^ {in1[20]});
 assign mul_34_17_n_982 = ~({in2[47]} ^ {in1[18]});
 assign mul_34_17_n_981 = ({in2[47]} ^ {in1[6]});
 assign mul_34_17_n_979 = ({in2[47]} ^ {in1[2]});
 assign mul_34_17_n_978 = ~({in2[47]} ^ {in1[26]});
 assign mul_34_17_n_977 = ({in2[47]} ^ {in1[4]});
 assign mul_34_17_n_976 = ({in2[47]} ^ {in1[29]});
 assign mul_34_17_n_974 = ~({in2[47]} ^ {in1[27]});
 assign mul_34_17_n_973 = ({in2[47]} ^ {in1[9]});
 assign mul_34_17_n_971 = ~({in2[47]} ^ {in1[22]});
 assign mul_34_17_n_969 = ({in2[47]} ^ {in1[3]});
 assign mul_34_17_n_968 = ({in2[47]} ^ {in1[35]});
 assign mul_34_17_n_967 = ({in2[49]} ^ {in1[1]});
 assign mul_34_17_n_965 = ~({in2[49]} ^ {in1[15]});
 assign mul_34_17_n_964 = ~({in2[49]} ^ {in1[21]});
 assign mul_34_17_n_962 = ~({in2[49]} ^ {in1[17]});
 assign mul_34_17_n_961 = ({in2[49]} ^ {in1[35]});
 assign mul_34_17_n_959 = ~({in2[49]} ^ {in1[28]});
 assign mul_34_17_n_958 = ~({in2[49]} ^ {in1[23]});
 assign mul_34_17_n_956 = ~({in2[49]} ^ {in1[19]});
 assign mul_34_17_n_955 = ({in2[25]} ^ {in1[36]});
 assign mul_34_17_n_953 = ~({in2[49]} ^ {in1[33]});
 assign mul_34_17_n_952 = ({in2[49]} ^ {in1[30]});
 assign mul_34_17_n_951 = ({in2[49]} ^ {in1[34]});
 assign mul_34_17_n_950 = ~({in2[49]} ^ {in1[12]});
 assign mul_34_17_n_949 = ~({in2[49]} ^ {in1[20]});
 assign mul_34_17_n_947 = ~({in2[49]} ^ {in1[14]});
 assign mul_34_17_n_946 = ({in2[49]} ^ {in1[4]});
 assign mul_34_17_n_945 = ({in2[49]} ^ {in1[3]});
 assign mul_34_17_n_944 = ({in2[49]} ^ {in1[25]});
 assign mul_34_17_n_943 = ({in2[49]} ^ {in1[18]});
 assign mul_34_17_n_941 = ~({in2[49]} ^ {in1[27]});
 assign mul_34_17_n_940 = ({in2[49]} ^ {in1[2]});
 assign mul_34_17_n_939 = ({in2[49]} ^ {in1[29]});
 assign mul_34_17_n_938 = ({in2[49]} ^ {in1[36]});
 assign mul_34_17_n_937 = ({in2[49]} ^ {in1[9]});
 assign mul_34_17_n_936 = ~({in2[61]} ^ {in1[17]});
 assign mul_34_17_n_934 = ~({in2[49]} ^ {in1[24]});
 assign mul_34_17_n_933 = ({in2[49]} ^ {in1[8]});
 assign mul_34_17_n_932 = ({in2[49]} ^ {in1[7]});
 assign mul_34_17_n_931 = ~({in2[49]} ^ {in1[11]});
 assign mul_34_17_n_929 = ~({in2[49]} ^ {in1[10]});
 assign mul_34_17_n_928 = ({in2[49]} ^ {in1[26]});
 assign mul_34_17_n_927 = ~({in2[49]} ^ {in1[22]});
 assign mul_34_17_n_926 = ~({in2[49]} ^ {in1[32]});
 assign mul_34_17_n_925 = ({in2[49]} ^ {in1[5]});
 assign mul_34_17_n_924 = ~({in2[49]} ^ {in1[16]});
 assign mul_34_17_n_923 = ({in2[49]} ^ {in1[6]});
 assign mul_34_17_n_921 = ~({in2[49]} ^ {in1[31]});
 assign mul_34_17_n_920 = ~({in2[49]} ^ {in1[13]});
 assign mul_34_17_n_918 = ~({in2[51]} ^ {in1[31]});
 assign mul_34_17_n_917 = ~({in2[51]} ^ {in1[20]});
 assign mul_34_17_n_916 = ({in2[51]} ^ {in1[3]});
 assign mul_34_17_n_915 = ({in2[51]} ^ {in1[4]});
 assign mul_34_17_n_913 = ({in2[51]} ^ {in1[12]});
 assign mul_34_17_n_912 = ({in2[51]} ^ {in1[33]});
 assign mul_34_17_n_911 = ({in2[51]} ^ {in1[34]});
 assign mul_34_17_n_910 = ({in2[51]} ^ {in1[1]});
 assign mul_34_17_n_909 = ({in2[51]} ^ {in1[5]});
 assign mul_34_17_n_908 = ~({in2[51]} ^ {in1[22]});
 assign mul_34_17_n_906 = ~({in2[51]} ^ {in1[18]});
 assign mul_34_17_n_905 = ({in2[51]} ^ {in1[28]});
 assign mul_34_17_n_904 = ~({in2[51]} ^ {in1[17]});
 assign mul_34_17_n_903 = ~({in2[25]} ^ {in1[38]});
 assign mul_34_17_n_902 = ~({in2[61]} ^ {in1[10]});
 assign mul_34_17_n_900 = ~({in2[51]} ^ {in1[19]});
 assign mul_34_17_n_899 = ~({in2[51]} ^ {in1[15]});
 assign mul_34_17_n_897 = ~({in2[51]} ^ {in1[10]});
 assign mul_34_17_n_896 = ~({in2[51]} ^ {in1[30]});
 assign mul_34_17_n_895 = ~({in2[51]} ^ {in1[13]});
 assign mul_34_17_n_894 = ~({in2[51]} ^ {in1[24]});
 assign mul_34_17_n_893 = ~({in2[51]} ^ {in1[8]});
 assign mul_34_17_n_892 = ({in2[51]} ^ {in1[2]});
 assign mul_34_17_n_891 = ~({in2[51]} ^ {in1[23]});
 assign mul_34_17_n_890 = ~({in2[51]} ^ {in1[25]});
 assign mul_34_17_n_889 = ({in2[51]} ^ {in1[11]});
 assign mul_34_17_n_888 = ({in2[51]} ^ {in1[6]});
 assign mul_34_17_n_887 = ~({in2[51]} ^ {in1[16]});
 assign mul_34_17_n_885 = ({in2[51]} ^ {in1[7]});
 assign mul_34_17_n_884 = ~({in2[51]} ^ {in1[9]});
 assign mul_34_17_n_882 = ~({in2[51]} ^ {in1[26]});
 assign mul_34_17_n_881 = ({in2[51]} ^ {in1[32]});
 assign mul_34_17_n_879 = ~({in2[51]} ^ {in1[29]});
 assign mul_34_17_n_878 = ~({in2[51]} ^ {in1[14]});
 assign mul_34_17_n_877 = ({in2[51]} ^ {in1[27]});
 assign mul_34_17_n_876 = ~({in2[51]} ^ {in1[21]});
 assign mul_34_17_n_874 = ({in2[53]} ^ {in1[2]});
 assign mul_34_17_n_872 = ~({in2[53]} ^ {in1[15]});
 assign mul_34_17_n_871 = ({in2[53]} ^ {in1[25]});
 assign mul_34_17_n_870 = ({in2[53]} ^ {in1[27]});
 assign mul_34_17_n_868 = ~({in2[53]} ^ {in1[1]});
 assign mul_34_17_n_867 = ~({in2[53]} ^ {in1[9]});
 assign mul_34_17_n_866 = ~({in2[25]} ^ {in1[50]});
 assign mul_34_17_n_865 = ({in2[53]} ^ {in1[26]});
 assign mul_34_17_n_864 = ~({in2[53]} ^ {in1[11]});
 assign mul_34_17_n_862 = ~({in2[53]} ^ {in1[28]});
 assign mul_34_17_n_861 = ({in2[53]} ^ {in1[14]});
 assign mul_34_17_n_859 = ~({in2[53]} ^ {in1[30]});
 assign mul_34_17_n_857 = ~({in2[53]} ^ {in1[6]});
 assign mul_34_17_n_856 = ({in2[53]} ^ {in1[31]});
 assign mul_34_17_n_855 = ({in2[53]} ^ {in1[5]});
 assign mul_34_17_n_854 = ({in2[53]} ^ {in1[32]});
 assign mul_34_17_n_853 = ({in2[53]} ^ {in1[23]});
 assign mul_34_17_n_852 = ({in2[53]} ^ {in1[22]});
 assign mul_34_17_n_851 = ~({in2[53]} ^ {in1[16]});
 assign mul_34_17_n_850 = ~({in2[53]} ^ {in1[18]});
 assign mul_34_17_n_849 = ~({in2[53]} ^ {in1[20]});
 assign mul_34_17_n_847 = ~({in2[53]} ^ {in1[21]});
 assign mul_34_17_n_846 = ~({in2[53]} ^ {in1[7]});
 assign mul_34_17_n_845 = ~({in2[53]} ^ {in1[19]});
 assign mul_34_17_n_844 = ~({in2[53]} ^ {in1[29]});
 assign mul_34_17_n_843 = ({in2[53]} ^ {in1[3]});
 assign mul_34_17_n_842 = ~({in2[61]} ^ {in1[6]});
 assign mul_34_17_n_840 = ~({in2[53]} ^ {in1[12]});
 assign mul_34_17_n_839 = ({in2[53]} ^ {in1[4]});
 assign mul_34_17_n_838 = ({in2[53]} ^ {in1[24]});
 assign mul_34_17_n_837 = ~({in2[53]} ^ {in1[10]});
 assign mul_34_17_n_836 = ~({in2[53]} ^ {in1[17]});
 assign mul_34_17_n_835 = ({in2[53]} ^ {in1[13]});
 assign mul_34_17_n_834 = ~({in2[53]} ^ {in1[8]});
 assign mul_34_17_n_833 = ~({in2[55]} ^ {in1[10]});
 assign mul_34_17_n_832 = ~({in2[55]} ^ {in1[23]});
 assign mul_34_17_n_831 = ~({in2[55]} ^ {in1[30]});
 assign mul_34_17_n_830 = ~({in2[55]} ^ {in1[11]});
 assign mul_34_17_n_829 = ~({in2[55]} ^ {in1[19]});
 assign mul_34_17_n_827 = ~({in2[25]} ^ {in1[41]});
 assign mul_34_17_n_826 = ~({in2[55]} ^ {in1[20]});
 assign mul_34_17_n_825 = ~({in2[55]} ^ {in1[2]});
 assign mul_34_17_n_824 = ~({in2[55]} ^ {in1[22]});
 assign mul_34_17_n_823 = ~({in2[55]} ^ {in1[16]});
 assign mul_34_17_n_822 = ~({in2[55]} ^ {in1[4]});
 assign mul_34_17_n_821 = ~({in2[55]} ^ {in1[9]});
 assign mul_34_17_n_820 = ~({in2[55]} ^ {in1[21]});
 assign mul_34_17_n_819 = ~({in2[55]} ^ {in1[14]});
 assign mul_34_17_n_818 = ~({in2[55]} ^ {in1[15]});
 assign mul_34_17_n_817 = ~({in2[55]} ^ {in1[28]});
 assign mul_34_17_n_816 = ~({in2[55]} ^ {in1[17]});
 assign mul_34_17_n_815 = ~({in2[55]} ^ {in1[25]});
 assign mul_34_17_n_814 = ~({in2[55]} ^ {in1[12]});
 assign mul_34_17_n_813 = ~({in2[55]} ^ {in1[13]});
 assign mul_34_17_n_812 = ~({in2[55]} ^ {in1[24]});
 assign mul_34_17_n_811 = ~({in2[55]} ^ {in1[26]});
 assign mul_34_17_n_810 = ~({in2[55]} ^ {in1[7]});
 assign mul_34_17_n_809 = ~({in2[55]} ^ {in1[18]});
 assign mul_34_17_n_808 = ~({in2[55]} ^ {in1[6]});
 assign mul_34_17_n_807 = ({in2[59]} ^ {in1[2]});
 assign mul_34_17_n_806 = ~({in2[55]} ^ {in1[29]});
 assign mul_34_17_n_805 = ~({in2[55]} ^ {in1[3]});
 assign mul_34_17_n_804 = ~({in2[55]} ^ {in1[8]});
 assign mul_34_17_n_803 = ~({in2[55]} ^ {in1[5]});
 assign mul_34_17_n_802 = ~({in2[55]} ^ {in1[1]});
 assign mul_34_17_n_801 = ~({in2[55]} ^ {in1[27]});
 assign mul_34_17_n_800 = ({in2[57]} ^ {in1[15]});
 assign mul_34_17_n_799 = ({in2[25]} ^ {in1[2]});
 assign mul_34_17_n_797 = ~({in2[57]} ^ {in1[10]});
 assign mul_34_17_n_796 = ({in2[57]} ^ {in1[23]});
 assign mul_34_17_n_795 = ({in2[57]} ^ {in1[26]});
 assign mul_34_17_n_794 = ({in2[57]} ^ {in1[20]});
 assign mul_34_17_n_793 = ~({in2[57]} ^ {in1[17]});
 assign mul_34_17_n_792 = ({in2[57]} ^ {in1[22]});
 assign mul_34_17_n_791 = ~({in2[57]} ^ {in1[13]});
 assign mul_34_17_n_790 = ({in2[57]} ^ {in1[8]});
 assign mul_34_17_n_789 = ({in2[57]} ^ {in1[21]});
 assign mul_34_17_n_788 = ({in2[57]} ^ {in1[28]});
 assign mul_34_17_n_786 = ~({in2[57]} ^ {in1[9]});
 assign mul_34_17_n_784 = ~({in2[57]} ^ {in1[24]});
 assign mul_34_17_n_782 = ~({in2[57]} ^ {in1[25]});
 assign mul_34_17_n_781 = ({in2[57]} ^ {in1[11]});
 assign mul_34_17_n_779 = ({in2[57]} ^ {in1[19]});
 assign mul_34_17_n_778 = ~({in2[57]} ^ {in1[18]});
 assign mul_34_17_n_777 = ({in2[57]} ^ {in1[27]});
 assign mul_34_17_n_775 = ~({in2[57]} ^ {in1[12]});
 assign mul_34_17_n_773 = ({in2[57]} ^ {in1[16]});
 assign mul_34_17_n_772 = ({in2[57]} ^ {in1[7]});
 assign mul_34_17_n_770 = ~({in2[57]} ^ {in1[6]});
 assign mul_34_17_n_769 = ~({in2[61]} ^ {in1[5]});
 assign mul_34_17_n_768 = ({in2[57]} ^ {in1[1]});
 assign mul_34_17_n_766 = ~({in2[57]} ^ {in1[14]});
 assign mul_34_17_n_765 = ({in2[57]} ^ {in1[4]});
 assign mul_34_17_n_763 = ~({in2[57]} ^ {in1[5]});
 assign mul_34_17_n_761 = ~({in2[57]} ^ {in1[3]});
 assign mul_34_17_n_759 = ~({in2[57]} ^ {in1[2]});
 assign mul_34_17_n_757 = ~({in2[59]} ^ {in1[23]});
 assign mul_34_17_n_755 = ~({in2[61]} ^ {in1[4]});
 assign mul_34_17_n_754 = ({in2[63]} ^ {in1[9]});
 assign mul_34_17_n_753 = ({in2[63]} ^ {in1[4]});
 assign mul_34_17_n_752 = ~({in2[61]} ^ {in1[21]});
 assign mul_34_17_n_751 = ({in2[63]} ^ {in1[5]});
 assign mul_34_17_n_750 = ({in2[59]} ^ {in1[21]});
 assign mul_34_17_n_748 = ~({in2[59]} ^ {in1[22]});
 assign mul_34_17_n_747 = ({in2[59]} ^ {in1[3]});
 assign mul_34_17_n_745 = ~({in2[63]} ^ {in1[13]});
 assign mul_34_17_n_744 = ({in2[59]} ^ {in1[6]});
 assign mul_34_17_n_743 = ({in2[59]} ^ {in1[20]});
 assign mul_34_17_n_741 = ~({in2[63]} ^ {in1[14]});
 assign mul_34_17_n_740 = ({in2[59]} ^ {in1[7]});
 assign mul_34_17_n_739 = ({in2[59]} ^ {in1[4]});
 assign mul_34_17_n_738 = ({in2[63]} ^ {in1[17]});
 assign mul_34_17_n_736 = ({in2[63]} ^ {in1[18]});
 assign mul_34_17_n_735 = ~({in2[59]} ^ {in1[17]});
 assign mul_34_17_n_734 = ({in2[63]} ^ {in1[2]});
 assign mul_34_17_n_733 = ~({in2[59]} ^ {in1[11]});
 assign mul_34_17_n_732 = ({in2[63]} ^ {in1[8]});
 assign mul_34_17_n_731 = ~({in2[61]} ^ {in1[12]});
 assign mul_34_17_n_730 = ~({in2[59]} ^ {in1[13]});
 assign mul_34_17_n_728 = ~({in2[63]} ^ {in1[20]});
 assign mul_34_17_n_727 = ~({in2[25]} ^ {in1[44]});
 assign mul_34_17_n_726 = ~({in2[61]} ^ {in1[1]});
 assign mul_34_17_n_725 = ~({in2[61]} ^ {in1[7]});
 assign mul_34_17_n_724 = ({in2[63]} ^ {in1[1]});
 assign mul_34_17_n_723 = ~({in2[61]} ^ {in1[8]});
 assign mul_34_17_n_722 = ~({in2[59]} ^ {in1[14]});
 assign mul_34_17_n_721 = ({in2[63]} ^ {in1[11]});
 assign mul_34_17_n_719 = ~({in2[63]} ^ {in1[7]});
 assign mul_34_17_n_718 = ({in2[59]} ^ {in1[19]});
 assign mul_34_17_n_716 = ~({in2[59]} ^ {in1[10]});
 assign mul_34_17_n_715 = ({in2[63]} ^ {in1[21]});
 assign mul_34_17_n_714 = ~({in2[59]} ^ {in1[15]});
 assign mul_34_17_n_713 = ~({in2[59]} ^ {in1[12]});
 assign mul_34_17_n_712 = ({in2[59]} ^ {in1[8]});
 assign mul_34_17_n_711 = ({in2[59]} ^ {in1[9]});
 assign mul_34_17_n_710 = ({in2[63]} ^ {in1[12]});
 assign mul_34_17_n_709 = ~({in2[61]} ^ {in1[23]});
 assign mul_34_17_n_708 = ~({in2[61]} ^ {in1[13]});
 assign mul_34_17_n_707 = ({in2[59]} ^ {in1[1]});
 assign mul_34_17_n_706 = ~({in2[61]} ^ {in1[3]});
 assign mul_34_17_n_705 = ({in2[63]} ^ {in1[15]});
 assign mul_34_17_n_704 = ~({in2[59]} ^ {in1[16]});
 assign mul_34_17_n_703 = ~({in2[61]} ^ {in1[2]});
 assign mul_34_17_n_702 = ~({in2[63]} ^ {in1[19]});
 assign mul_34_17_n_701 = ~({in2[61]} ^ {in1[18]});
 assign mul_34_17_n_700 = ~({in2[61]} ^ {in1[9]});
 assign mul_34_17_n_699 = ({in2[63]} ^ {in1[3]});
 assign mul_34_17_n_698 = ~({in2[61]} ^ {in1[15]});
 assign mul_34_17_n_697 = ~({in2[61]} ^ {in1[14]});
 assign mul_34_17_n_696 = ~({in2[61]} ^ {in1[11]});
 assign mul_34_17_n_695 = ({in2[59]} ^ {in1[5]});
 assign mul_34_17_n_694 = ~({in2[61]} ^ {in1[19]});
 assign mul_34_17_n_693 = ({in2[63]} ^ {in1[22]});
 assign mul_34_17_n_692 = ~({in2[61]} ^ {in1[16]});
 assign mul_34_17_n_691 = ({in2[61]} ^ {in2[62]});
 assign mul_34_17_n_689 = ({in2[59]} ^ {in2[60]});
 assign mul_34_17_n_687 = ({in2[57]} ^ {in2[58]});
 assign mul_34_17_n_685 = ({in2[55]} ^ {in2[56]});
 assign mul_34_17_n_683 = ({in2[53]} ^ {in2[54]});
 assign mul_34_17_n_681 = ({in2[51]} ^ {in2[52]});
 assign mul_34_17_n_679 = ({in2[49]} ^ {in2[50]});
 assign mul_34_17_n_677 = ({in2[47]} ^ {in2[48]});
 assign mul_34_17_n_675 = ({in2[45]} ^ {in2[46]});
 assign mul_34_17_n_673 = ({in2[43]} ^ {in2[44]});
 assign mul_34_17_n_671 = ({in2[41]} ^ {in2[42]});
 assign mul_34_17_n_669 = ({in2[39]} ^ {in2[40]});
 assign mul_34_17_n_667 = ({in2[37]} ^ {in2[38]});
 assign mul_34_17_n_665 = ({in2[35]} ^ {in2[36]});
 assign mul_34_17_n_663 = ({in2[33]} ^ {in2[34]});
 assign mul_34_17_n_661 = ({in2[31]} ^ {in2[32]});
 assign mul_34_17_n_659 = ({in2[29]} ^ {in2[30]});
 assign mul_34_17_n_657 = ({in2[27]} ^ {in2[28]});
 assign mul_34_17_n_655 = ({in2[25]} ^ {in2[26]});
 assign mul_34_17_n_571 = ~({in2[56]} | {in1[0]});
 assign mul_34_17_n_570 = ~({in2[56]} & {in1[0]});
 assign mul_34_17_n_569 = ~({in2[54]} & {in1[0]});
 assign mul_34_17_n_568 = ~({in2[50]} | {in1[0]});
 assign mul_34_17_n_567 = ~({in2[28]} | {in1[0]});
 assign mul_34_17_n_566 = ~({in2[48]} | {in1[0]});
 assign mul_34_17_n_565 = ~({in2[26]} & {in1[0]});
 assign mul_34_17_n_564 = ~({in2[32]} | {in1[0]});
 assign mul_34_17_n_563 = ~({in2[12]} & {in1[0]});
 assign mul_34_17_n_562 = ~({in2[42]} | {in1[0]});
 assign mul_34_17_n_561 = ~({in2[18]} & {in1[0]});
 assign mul_34_17_n_560 = ~({in2[26]} | {in1[0]});
 assign mul_34_17_n_559 = ~({in2[12]} | {in1[0]});
 assign mul_34_17_n_558 = ~({in2[22]} & {in1[0]});
 assign mul_34_17_n_557 = ~({in2[2]} & {in1[0]});
 assign mul_34_17_n_556 = ~({in2[58]} & {in1[0]});
 assign mul_34_17_n_555 = ~({in2[22]} | {in1[0]});
 assign mul_34_17_n_554 = ~({in2[34]} & {in1[0]});
 assign mul_34_17_n_553 = ~({in2[40]} & {in1[0]});
 assign mul_34_17_n_552 = ~({in2[34]} | {in1[0]});
 assign mul_34_17_n_551 = ~({in2[54]} | {in1[0]});
 assign mul_34_17_n_550 = ~({in2[52]} & {in1[0]});
 assign mul_34_17_n_549 = ~({in2[10]} | {in1[0]});
 assign mul_34_17_n_548 = ~({in2[38]} | {in1[0]});
 assign mul_34_17_n_547 = ~({in2[20]} | {in1[0]});
 assign mul_34_17_n_546 = ~({in2[60]} & {in1[0]});
 assign mul_34_17_n_545 = ~({in2[50]} & {in1[0]});
 assign mul_34_17_n_544 = ~({in2[30]} | {in1[0]});
 assign mul_34_17_n_543 = ~({in2[44]} & {in1[0]});
 assign mul_34_17_n_542 = ~({in2[24]} | {in1[0]});
 assign mul_34_17_n_541 = ~({in2[28]} & {in1[0]});
 assign mul_34_17_n_540 = ~({in2[58]} | {in1[0]});
 assign mul_34_17_n_539 = ~({in2[32]} & {in1[0]});
 assign mul_34_17_n_538 = ~({in2[52]} | {in1[0]});
 assign mul_34_17_n_537 = ~({in2[10]} & {in1[0]});
 assign mul_34_17_n_536 = ~({in2[8]} | {in1[0]});
 assign mul_34_17_n_535 = ~({in2[38]} & {in1[0]});
 assign mul_34_17_n_534 = ~({in2[24]} & {in1[0]});
 assign mul_34_17_n_533 = ~({in2[48]} & {in1[0]});
 assign mul_34_17_n_532 = ~({in2[16]} | {in1[0]});
 assign mul_34_17_n_531 = ~({in2[2]} | {in1[0]});
 assign mul_34_17_n_518 = ~mul_34_17_n_517;
 assign mul_34_17_n_515 = ~({in2[53]} & {in1[0]});
 assign mul_34_17_n_514 = ~({in2[4]} & {in1[0]});
 assign mul_34_17_n_513 = ~({in2[46]} | {in1[0]});
 assign mul_34_17_n_512 = ~({in2[36]} | {in1[0]});
 assign mul_34_17_n_511 = ~({in2[18]} | {in1[0]});
 assign mul_34_17_n_510 = ~({in2[16]} & {in1[0]});
 assign mul_34_17_n_509 = ~({in2[60]} | {in1[0]});
 assign mul_34_17_n_508 = ~({in2[14]} | {in1[0]});
 assign mul_34_17_n_507 = ~({in2[42]} & {in1[0]});
 assign mul_34_17_n_506 = ~({in2[20]} & {in1[0]});
 assign mul_34_17_n_505 = ~({in2[30]} & {in1[0]});
 assign mul_34_17_n_504 = ~({in2[62]} | {in1[0]});
 assign mul_34_17_n_503 = ~({in2[8]} & {in1[0]});
 assign mul_34_17_n_502 = ~({in2[46]} & {in1[0]});
 assign mul_34_17_n_501 = ~({in2[6]} & {in1[0]});
 assign mul_34_17_n_500 = ~({in2[36]} & {in1[0]});
 assign mul_34_17_n_499 = ~({in2[62]} & {in1[0]});
 assign mul_34_17_n_498 = ~({in2[14]} & {in1[0]});
 assign mul_34_17_n_497 = ~({in2[40]} | {in1[0]});
 assign mul_34_17_n_496 = ~({in2[44]} | {in1[0]});
 assign mul_34_17_n_495 = ~({in2[6]} | {in1[0]});
 assign mul_34_17_n_530 = ~(mul_34_17_n_426 & {in2[19]});
 assign mul_34_17_n_494 = ~({in1[63]} | mul_34_17_n_416);
 assign mul_34_17_n_493 = ~({in2[21]} | mul_34_17_n_426);
 assign mul_34_17_n_529 = ~({in1[63]} | mul_34_17_n_417);
 assign mul_34_17_n_492 = ~({in2[15]} | mul_34_17_n_426);
 assign mul_34_17_n_528 = ~({in1[63]} | mul_34_17_n_418);
 assign mul_34_17_n_527 = ~({in2[11]} | mul_34_17_n_426);
 assign mul_34_17_n_526 = ~({in1[63]} | mul_34_17_n_394);
 assign mul_34_17_n_491 = ~(mul_34_17_n_396 & {in1[63]});
 assign mul_34_17_n_525 = ~({in2[9]} | mul_34_17_n_426);
 assign mul_34_17_n_524 = ~({in1[63]} | mul_34_17_n_415);
 assign mul_34_17_n_490 = ~(mul_34_17_n_426 & {in2[7]});
 assign mul_34_17_n_523 = ~({in2[13]} | mul_34_17_n_426);
 assign mul_34_17_n_489 = ~({in2[3]} | mul_34_17_n_426);
 assign mul_34_17_n_488 = ~({in1[63]} | mul_34_17_n_413);
 assign mul_34_17_n_522 = ~({in2[17]} | mul_34_17_n_426);
 assign mul_34_17_n_487 = ~({in1[63]} | mul_34_17_n_393);
 assign mul_34_17_n_521 = ~(mul_34_17_n_426 & {in2[5]});
 assign mul_34_17_n_520 = ~(mul_34_17_n_395 & {in1[63]});
 assign mul_34_17_n_519 = ~(mul_34_17_n_412 & {in1[63]});
 assign mul_34_17_n_486 = ~({in1[63]} | mul_34_17_n_397);
 assign mul_34_17_n_485 = ~({in2[1]} | mul_34_17_n_426);
 assign mul_34_17_n_484 = ~({in2[63]} | {in1[0]});
 assign mul_34_17_n_483 = ~({in2[63]} & {in1[0]});
 assign mul_34_17_n_482 = ~({in2[59]} | {in1[0]});
 assign mul_34_17_n_481 = ~({in2[59]} & {in1[0]});
 assign mul_34_17_n_480 = ~({in2[57]} & {in1[0]});
 assign mul_34_17_n_479 = ~({in2[57]} | {in1[0]});
 assign mul_34_17_n_478 = ~({in2[19]} & {in1[0]});
 assign mul_34_17_n_477 = ~({in2[53]} | {in1[0]});
 assign mul_34_17_n_476 = ~({in2[4]} | {in1[0]});
 assign mul_34_17_n_475 = ~({in2[51]} | {in1[0]});
 assign mul_34_17_n_474 = ~({in2[51]} & {in1[0]});
 assign mul_34_17_n_473 = ~({in2[49]} & {in1[0]});
 assign mul_34_17_n_472 = ~({in2[49]} | {in1[0]});
 assign mul_34_17_n_471 = ~({in2[47]} | {in1[0]});
 assign mul_34_17_n_470 = ~({in2[47]} & {in1[0]});
 assign mul_34_17_n_469 = ~({in2[45]} | {in1[0]});
 assign mul_34_17_n_468 = ~({in2[45]} & {in1[0]});
 assign mul_34_17_n_467 = ~({in2[43]} | {in1[0]});
 assign mul_34_17_n_466 = ~({in2[43]} & {in1[0]});
 assign mul_34_17_n_465 = ~({in2[41]} & {in1[0]});
 assign mul_34_17_n_464 = ~({in2[41]} | {in1[0]});
 assign mul_34_17_n_463 = ~({in2[39]} | {in1[0]});
 assign mul_34_17_n_462 = ~({in2[39]} & {in1[0]});
 assign mul_34_17_n_461 = ~({in2[37]} | {in1[0]});
 assign mul_34_17_n_460 = ~({in2[37]} & {in1[0]});
 assign mul_34_17_n_459 = ~({in2[35]} & {in1[0]});
 assign mul_34_17_n_458 = ~({in2[35]} | {in1[0]});
 assign mul_34_17_n_457 = ~({in2[33]} & {in1[0]});
 assign mul_34_17_n_456 = ~({in2[33]} | {in1[0]});
 assign mul_34_17_n_455 = ~({in2[23]} | {in1[0]});
 assign mul_34_17_n_454 = ~({in2[31]} & {in1[0]});
 assign mul_34_17_n_453 = ~({in2[31]} | {in1[0]});
 assign mul_34_17_n_452 = ~({in2[29]} & {in1[0]});
 assign mul_34_17_n_451 = ~({in2[29]} | {in1[0]});
 assign mul_34_17_n_450 = ~({in2[27]} | {in1[0]});
 assign mul_34_17_n_449 = ~({in2[27]} & {in1[0]});
 assign mul_34_17_n_448 = ~({in2[25]} & {in1[0]});
 assign mul_34_17_n_447 = ~({in2[25]} | {in1[0]});
 assign mul_34_17_n_446 = ~({in2[3]} | {in1[0]});
 assign mul_34_17_n_445 = ~({in2[21]} & {in1[0]});
 assign mul_34_17_n_444 = ~({in2[11]} & {in1[0]});
 assign mul_34_17_n_443 = ~({in2[19]} | {in1[0]});
 assign mul_34_17_n_442 = ~({in2[7]} | {in1[0]});
 assign mul_34_17_n_441 = ~({in2[11]} | {in1[0]});
 assign mul_34_17_n_440 = ~({in2[9]} | {in1[0]});
 assign mul_34_17_n_439 = ~({in2[21]} | {in1[0]});
 assign mul_34_17_n_438 = ~({in2[17]} | {in1[0]});
 assign mul_34_17_n_437 = ~({in2[3]} & {in1[0]});
 assign mul_34_17_n_436 = ~({in2[7]} & {in1[0]});
 assign mul_34_17_n_435 = ~({in2[23]} & {in1[0]});
 assign mul_34_17_n_434 = ~({in2[17]} & {in1[0]});
 assign mul_34_17_n_433 = ~({in2[13]} & {in1[0]});
 assign mul_34_17_n_432 = ~({in2[15]} & {in1[0]});
 assign mul_34_17_n_431 = ~({in2[13]} | {in1[0]});
 assign mul_34_17_n_430 = ~({in2[5]} & {in1[0]});
 assign mul_34_17_n_429 = ~({in2[15]} | {in1[0]});
 assign mul_34_17_n_428 = ~({in2[9]} & {in1[0]});
 assign mul_34_17_n_427 = ~({in2[5]} | {in1[0]});
 assign mul_34_17_n_517 = ~({in2[0]} & {in1[0]});
 assign mul_34_17_n_516 = ~({in2[0]} | mul_34_17_n_397);
 assign mul_34_17_n_426 = ~{in1[63]};
 assign mul_34_17_n_425 = ~{in2[63]};
 assign mul_34_17_n_424 = ~{in2[61]};
 assign mul_34_17_n_423 = ~{in2[57]};
 assign mul_34_17_n_422 = ~{in2[55]};
 assign mul_34_17_n_421 = ~{in2[49]};
 assign mul_34_17_n_420 = ~{in2[45]};
 assign mul_34_17_n_419 = ~{in2[37]};
 assign mul_34_17_n_418 = ~{in2[11]};
 assign mul_34_17_n_417 = ~{in2[9]};
 assign mul_34_17_n_416 = ~{in2[21]};
 assign mul_34_17_n_415 = ~{in2[17]};
 assign mul_34_17_n_414 = ~{in2[23]};
 assign mul_34_17_n_413 = ~{in2[3]};
 assign mul_34_17_n_412 = ~{in2[5]};
 assign mul_34_17_n_411 = ~{in1[0]};
 assign mul_34_17_n_410 = ~{in2[59]};
 assign mul_34_17_n_409 = ~{in2[53]};
 assign mul_34_17_n_408 = ~{in2[51]};
 assign mul_34_17_n_407 = ~{in2[47]};
 assign mul_34_17_n_406 = ~{in2[43]};
 assign mul_34_17_n_405 = ~{in2[41]};
 assign mul_34_17_n_404 = ~{in2[39]};
 assign mul_34_17_n_403 = ~{in2[35]};
 assign mul_34_17_n_402 = ~{in2[33]};
 assign mul_34_17_n_401 = ~{in2[31]};
 assign mul_34_17_n_400 = ~{in2[29]};
 assign mul_34_17_n_399 = ~{in2[27]};
 assign mul_34_17_n_398 = ~{in2[25]};
 assign mul_34_17_n_397 = ~{in2[1]};
 assign mul_34_17_n_396 = ~{in2[7]};
 assign mul_34_17_n_395 = ~{in2[19]};
 assign mul_34_17_n_394 = ~{in2[13]};
 assign mul_34_17_n_393 = ~{in2[15]};
 assign mul_34_17_n_390 = ((mul_34_17_n_2832 & mul_34_17_n_4288) | ((mul_34_17_n_2832 & mul_34_17_n_2718)
    | (mul_34_17_n_2718 & mul_34_17_n_4288)));
 assign mul_34_17_n_389 = (mul_34_17_n_5517 ^ mul_34_17_n_5509);
 assign mul_34_17_n_388 = ~(mul_34_17_n_6342 ^ mul_34_17_n_6341);
 assign mul_34_17_n_387 = (mul_34_17_n_6471 ^ mul_34_17_n_2);
 assign mul_34_17_n_386 = ~(mul_34_17_n_6785 ^ mul_34_17_n_5508);
 assign mul_34_17_n_385 = ~(mul_34_17_n_6338 ^ mul_34_17_n_5920);
 assign mul_34_17_n_384 = ~(mul_34_17_n_7306 ^ mul_34_17_n_30);
 assign mul_34_17_n_383 = (mul_34_17_n_135 ^ mul_34_17_n_146);
 assign mul_34_17_n_382 = (mul_34_17_n_6483 ^ mul_34_17_n_6525);
 assign mul_34_17_n_381 = (mul_34_17_n_6481 ^ mul_34_17_n_6501);
 assign mul_34_17_n_380 = ~(mul_34_17_n_7669 ^ mul_34_17_n_7439);
 assign mul_34_17_n_379 = ~(mul_34_17_n_6538 ^ mul_34_17_n_6541);
 assign mul_34_17_n_378 = (mul_34_17_n_7761 ^ mul_34_17_n_6776);
 assign mul_34_17_n_377 = (mul_34_17_n_7065 ^ mul_34_17_n_7049);
 assign mul_34_17_n_376 = (mul_34_17_n_6243 ^ mul_34_17_n_6240);
 assign mul_34_17_n_375 = ~(mul_34_17_n_7061 ^ mul_34_17_n_6462);
 assign mul_34_17_n_374 = ~(mul_34_17_n_7678 ^ mul_34_17_n_6894);
 assign mul_34_17_n_373 = (mul_34_17_n_7100 ^ mul_34_17_n_7118);
 assign mul_34_17_n_372 = (mul_34_17_n_7411 ^ mul_34_17_n_7429);
 assign mul_34_17_n_371 = (mul_34_17_n_7839 ^ mul_34_17_n_7846);
 assign mul_34_17_n_370 = ~(mul_34_17_n_7852 ^ mul_34_17_n_7981);
 assign mul_34_17_n_369 = ~(mul_34_17_n_6790 ^ mul_34_17_n_5107);
 assign mul_34_17_n_368 = ~(mul_34_17_n_7499 ^ mul_34_17_n_7494);
 assign mul_34_17_n_367 = ~(mul_34_17_n_11489 ^ mul_34_17_n_7410);
 assign mul_34_17_n_366 = ~(mul_34_17_n_11416 ^ mul_34_17_n_7854);
 assign mul_34_17_n_365 = (mul_34_17_n_11408 ^ mul_34_17_n_11412);
 assign mul_34_17_n_364 = ~(mul_34_17_n_8223 ^ mul_34_17_n_7668);
 assign mul_34_17_n_363 = ~(mul_34_17_n_8141 ^ mul_34_17_n_7762);
 assign mul_34_17_n_362 = ~(mul_34_17_n_8767 ^ mul_34_17_n_8486);
 assign mul_34_17_n_361 = ~(mul_34_17_n_8918 ^ mul_34_17_n_8731);
 assign mul_34_17_n_360 = ~(mul_34_17_n_8611 ^ mul_34_17_n_8593);
 assign mul_34_17_n_359 = (mul_34_17_n_8733 ^ mul_34_17_n_8493);
 assign mul_34_17_n_358 = ~(mul_34_17_n_9002 ^ mul_34_17_n_8645);
 assign mul_34_17_n_357 = ~(mul_34_17_n_9263 ^ mul_34_17_n_8829);
 assign mul_34_17_n_356 = (mul_34_17_n_9261 ^ mul_34_17_n_8982);
 assign mul_34_17_n_355 = ~(mul_34_17_n_9273 ^ mul_34_17_n_8726);
 assign mul_34_17_n_354 = ~(mul_34_17_n_9327 ^ mul_34_17_n_9462);
 assign mul_34_17_n_353 = (mul_34_17_n_9326 ^ mul_34_17_n_9411);
 assign mul_34_17_n_352 = ~(mul_34_17_n_9541 ^ mul_34_17_n_9088);
 assign mul_34_17_n_351 = ((mul_34_17_n_9265 & mul_34_17_n_9487) | ((mul_34_17_n_9265 & mul_34_17_n_9464)
    | (mul_34_17_n_9464 & mul_34_17_n_9487)));
 assign mul_34_17_n_350 = ~(mul_34_17_n_283 ^ mul_34_17_n_9480);
 assign mul_34_17_n_348 = ~mul_34_17_n_349;
 assign mul_34_17_n_349 = ~(mul_34_17_n_10082 | mul_34_17_n_10248);
 assign mul_34_17_n_346 = ~mul_34_17_n_347;
 assign mul_34_17_n_347 = ~(mul_34_17_n_9995 & mul_34_17_n_10214);
 assign mul_34_17_n_344 = ~mul_34_17_n_345;
 assign mul_34_17_n_345 = ~(mul_34_17_n_10094 | mul_34_17_n_10165);
 assign mul_34_17_n_342 = ~mul_34_17_n_343;
 assign mul_34_17_n_343 = ~(mul_34_17_n_10161 & mul_34_17_n_10164);
 assign mul_34_17_n_340 = ~mul_34_17_n_341;
 assign mul_34_17_n_341 = ~(mul_34_17_n_10103 & mul_34_17_n_9932);
 assign mul_34_17_n_339 = (mul_34_17_n_10136 ^ mul_34_17_n_10098);
 assign mul_34_17_n_338 = (mul_34_17_n_10138 ^ mul_34_17_n_10097);
 assign mul_34_17_n_337 = (mul_34_17_n_10191 ^ mul_34_17_n_10083);
 assign mul_34_17_n_335 = ~mul_34_17_n_336;
 assign mul_34_17_n_336 = ~(mul_34_17_n_9811 | mul_34_17_n_10028);
 assign mul_34_17_n_333 = ~mul_34_17_n_334;
 assign mul_34_17_n_334 = ~(mul_34_17_n_9973 | mul_34_17_n_9825);
 assign mul_34_17_n_332 = (mul_34_17_n_9960 ^ mul_34_17_n_9897);
 assign mul_34_17_n_330 = ~mul_34_17_n_331;
 assign mul_34_17_n_331 = ~(mul_34_17_n_9729 | mul_34_17_n_303);
 assign mul_34_17_n_328 = ~mul_34_17_n_329;
 assign mul_34_17_n_329 = ~(mul_34_17_n_9914 & mul_34_17_n_11282);
 assign mul_34_17_n_327 = (mul_34_17_n_9909 ^ mul_34_17_n_10064);
 assign mul_34_17_n_325 = ~mul_34_17_n_326;
 assign mul_34_17_n_326 = ~(mul_34_17_n_318 | mul_34_17_n_9907);
 assign mul_34_17_n_323 = ~mul_34_17_n_324;
 assign mul_34_17_n_324 = ~(mul_34_17_n_9877 & mul_34_17_n_9561);
 assign mul_34_17_n_322 = (mul_34_17_n_9935 ^ mul_34_17_n_9830);
 assign mul_34_17_n_321 = (mul_34_17_n_9824 ^ mul_34_17_n_9823);
 assign mul_34_17_n_319 = ~mul_34_17_n_320;
 assign mul_34_17_n_320 = ~(mul_34_17_n_9678 | mul_34_17_n_294);
 assign mul_34_17_n_318 = (mul_34_17_n_9691 ^ mul_34_17_n_9733);
 assign mul_34_17_n_317 = (mul_34_17_n_9692 ^ mul_34_17_n_9731);
 assign mul_34_17_n_315 = ~mul_34_17_n_316;
 assign mul_34_17_n_316 = ~(mul_34_17_n_9530 | mul_34_17_n_9664);
 assign mul_34_17_n_313 = ~mul_34_17_n_314;
 assign mul_34_17_n_314 = ~(mul_34_17_n_9369 | mul_34_17_n_9627);
 assign mul_34_17_n_311 = ~mul_34_17_n_312;
 assign mul_34_17_n_312 = ~(mul_34_17_n_9199 | mul_34_17_n_9617);
 assign mul_34_17_n_309 = ~mul_34_17_n_310;
 assign mul_34_17_n_310 = ~(mul_34_17_n_9596 | mul_34_17_n_9595);
 assign mul_34_17_n_308 = (mul_34_17_n_9536 ^ mul_34_17_n_9527);
 assign mul_34_17_n_306 = (mul_34_17_n_9365 ^ mul_34_17_n_9501);
 assign mul_34_17_n_305 = ~mul_34_17_n_391;
 assign mul_34_17_n_391 = ~(mul_34_17_n_9374 | mul_34_17_n_9499);
 assign mul_34_17_n_304 = (mul_34_17_n_9262 ^ mul_34_17_n_9474);
 assign mul_34_17_n_303 = (mul_34_17_n_9425 ^ mul_34_17_n_9698);
 assign mul_34_17_n_301 = ~mul_34_17_n_302;
 assign mul_34_17_n_302 = ~(mul_34_17_n_9376 | mul_34_17_n_9304);
 assign mul_34_17_n_300 = (mul_34_17_n_9745 ^ mul_34_17_n_9359);
 assign mul_34_17_n_299 = (mul_34_17_n_8985 ^ mul_34_17_n_9355);
 assign mul_34_17_n_294 = (mul_34_17_n_9453 ^ mul_34_17_n_9205);
 assign mul_34_17_n_292 = (mul_34_17_n_9449 ^ mul_34_17_n_9184);
 assign mul_34_17_n_291 = (mul_34_17_n_9628 ^ mul_34_17_n_9159);
 assign mul_34_17_n_290 = (mul_34_17_n_9061 ^ mul_34_17_n_9129);
 assign mul_34_17_n_287 = (mul_34_17_n_8995 ^ mul_34_17_n_9310);
 assign mul_34_17_n_286 = (mul_34_17_n_9063 ^ mul_34_17_n_8935);
 assign mul_34_17_n_285 = (mul_34_17_n_8963 ^ mul_34_17_n_8875);
 assign mul_34_17_n_284 = (mul_34_17_n_8870 ^ mul_34_17_n_8333);
 assign mul_34_17_n_283 = (mul_34_17_n_9059 ^ mul_34_17_n_8786);
 assign mul_34_17_n_282 = (mul_34_17_n_8883 ^ mul_34_17_n_8780);
 assign mul_34_17_n_281 = (mul_34_17_n_9058 ^ mul_34_17_n_8756);
 assign mul_34_17_n_280 = (mul_34_17_n_9064 ^ mul_34_17_n_8678);
 assign mul_34_17_n_279 = (mul_34_17_n_9060 ^ mul_34_17_n_11362);
 assign mul_34_17_n_278 = (mul_34_17_n_8966 ^ mul_34_17_n_8666);
 assign mul_34_17_n_277 = (mul_34_17_n_8968 ^ mul_34_17_n_8663);
 assign mul_34_17_n_276 = (mul_34_17_n_284 ^ mul_34_17_n_8612);
 assign mul_34_17_n_275 = (mul_34_17_n_8583 ^ mul_34_17_n_8567);
 assign mul_34_17_n_274 = (mul_34_17_n_8967 ^ mul_34_17_n_8566);
 assign mul_34_17_n_273 = (mul_34_17_n_8437 ^ mul_34_17_n_8565);
 assign mul_34_17_n_272 = (mul_34_17_n_8817 ^ mul_34_17_n_8560);
 assign mul_34_17_n_271 = (mul_34_17_n_8824 ^ mul_34_17_n_8558);
 assign mul_34_17_n_270 = (mul_34_17_n_8884 ^ mul_34_17_n_8551);
 assign mul_34_17_n_269 = (mul_34_17_n_8548 ^ mul_34_17_n_8226);
 assign mul_34_17_n_268 = (mul_34_17_n_8888 ^ mul_34_17_n_8536);
 assign mul_34_17_n_267 = (mul_34_17_n_8893 ^ mul_34_17_n_8513);
 assign mul_34_17_n_266 = (mul_34_17_n_8285 ^ mul_34_17_n_8412);
 assign mul_34_17_n_265 = (mul_34_17_n_8937 ^ mul_34_17_n_8356);
 assign mul_34_17_n_264 = (mul_34_17_n_8298 ^ mul_34_17_n_8267);
 assign mul_34_17_n_263 = (mul_34_17_n_8295 ^ mul_34_17_n_8264);
 assign mul_34_17_n_261 = ~mul_34_17_n_262;
 assign mul_34_17_n_262 = ~(mul_34_17_n_7998 & mul_34_17_n_8253);
 assign mul_34_17_n_260 = (mul_34_17_n_8811 ^ mul_34_17_n_8246);
 assign mul_34_17_n_259 = (mul_34_17_n_8283 ^ mul_34_17_n_8148);
 assign mul_34_17_n_257 = (mul_34_17_n_8079 ^ mul_34_17_n_7793);
 assign mul_34_17_n_256 = (mul_34_17_n_8087 ^ mul_34_17_n_7791);
 assign mul_34_17_n_255 = (mul_34_17_n_8197 ^ mul_34_17_n_11483);
 assign mul_34_17_n_254 = (mul_34_17_n_8440 ^ mul_34_17_n_7749);
 assign mul_34_17_n_253 = (mul_34_17_n_8063 ^ mul_34_17_n_7735);
 assign mul_34_17_n_251 = (mul_34_17_n_8194 ^ mul_34_17_n_7695);
 assign mul_34_17_n_249 = ~mul_34_17_n_250;
 assign mul_34_17_n_250 = ~(mul_34_17_n_7598 & mul_34_17_n_6776);
 assign mul_34_17_n_247 = (mul_34_17_n_7809 ^ mul_34_17_n_11494);
 assign mul_34_17_n_246 = (mul_34_17_n_8084 ^ mul_34_17_n_7568);
 assign mul_34_17_n_244 = (mul_34_17_n_8438 ^ mul_34_17_n_7541);
 assign mul_34_17_n_242 = ~mul_34_17_n_243;
 assign mul_34_17_n_243 = ~(mul_34_17_n_369 & mul_34_17_n_7066);
 assign mul_34_17_n_241 = (mul_34_17_n_239 ^ mul_34_17_n_11504);
 assign mul_34_17_n_240 = (mul_34_17_n_8443 ^ mul_34_17_n_7476);
 assign mul_34_17_n_239 = (mul_34_17_n_211 ^ mul_34_17_n_7464);
 assign mul_34_17_n_237 = ~mul_34_17_n_238;
 assign mul_34_17_n_238 = ~(mul_34_17_n_7459 | mul_34_17_n_7436);
 assign mul_34_17_n_236 = (mul_34_17_n_11394 ^ (mul_34_17_n_8036 ^ (mul_34_17_n_8132 ^ mul_34_17_n_7437)));
 assign mul_34_17_n_235 = (mul_34_17_n_8135 ^ mul_34_17_n_7423);
 assign mul_34_17_n_234 = (mul_34_17_n_8041 ^ mul_34_17_n_166);
 assign mul_34_17_n_233 = (mul_34_17_n_7951 ^ mul_34_17_n_7380);
 assign mul_34_17_n_232 = (mul_34_17_n_7178 ^ mul_34_17_n_7361);
 assign mul_34_17_n_231 = (mul_34_17_n_7952 ^ mul_34_17_n_7335);
 assign mul_34_17_n_230 = (mul_34_17_n_8287 ^ mul_34_17_n_7312);
 assign mul_34_17_n_229 = (mul_34_17_n_6953 ^ mul_34_17_n_7141);
 assign mul_34_17_n_228 = (mul_34_17_n_7182 ^ mul_34_17_n_7139);
 assign mul_34_17_n_227 = (mul_34_17_n_6952 ^ mul_34_17_n_7132);
 assign mul_34_17_n_226 = (mul_34_17_n_7817 ^ mul_34_17_n_7098);
 assign mul_34_17_n_225 = ((mul_34_17_n_149 & mul_34_17_n_7061) | ((mul_34_17_n_149 & mul_34_17_n_6462)
    | (mul_34_17_n_6462 & mul_34_17_n_7061)));
 assign mul_34_17_n_224 = (mul_34_17_n_6958 ^ mul_34_17_n_6923);
 assign mul_34_17_n_223 = ~((mul_34_17_n_7273 & ~mul_34_17_n_107) | (mul_34_17_n_7230 & mul_34_17_n_107));
 assign mul_34_17_n_221 = (mul_34_17_n_7172 ^ mul_34_17_n_53);
 assign mul_34_17_n_219 = (mul_34_17_n_7180 ^ (mul_34_17_n_6625 ^ (mul_34_17_n_7386 ^ mul_34_17_n_5912)));
 assign mul_34_17_n_218 = (mul_34_17_n_7168 ^ mul_34_17_n_6591);
 assign mul_34_17_n_215 = (mul_34_17_n_6661 ^ (mul_34_17_n_28 ^ (mul_34_17_n_5492 ^ mul_34_17_n_4429)));
 assign mul_34_17_n_213 = ~(mul_34_17_n_6384 ^ (mul_34_17_n_6348 ^ (mul_34_17_n_5495 ^ mul_34_17_n_3817)));
 assign mul_34_17_n_211 = ~((mul_34_17_n_7038 & ~mul_34_17_n_11) | (mul_34_17_n_7245 & mul_34_17_n_11));
 assign mul_34_17_n_209 = ~mul_34_17_n_210;
 assign mul_34_17_n_210 = ~(mul_34_17_n_6298 & mul_34_17_n_5521);
 assign mul_34_17_n_207 = (mul_34_17_n_7094 ^ mul_34_17_n_6161);
 assign mul_34_17_n_206 = (mul_34_17_n_7111 ^ mul_34_17_n_26);
 assign mul_34_17_n_204 = ~mul_34_17_n_205;
 assign mul_34_17_n_205 = ~(mul_34_17_n_6115 & mul_34_17_n_2867);
 assign mul_34_17_n_202 = ~mul_34_17_n_203;
 assign mul_34_17_n_203 = ((mul_34_17_n_5611 & mul_34_17_n_6112) | ((mul_34_17_n_5611 & mul_34_17_n_6004)
    | (mul_34_17_n_6004 & mul_34_17_n_6112)));
 assign mul_34_17_n_201 = (mul_34_17_n_6944 ^ mul_34_17_n_6111);
 assign mul_34_17_n_199 = ~mul_34_17_n_200;
 assign mul_34_17_n_200 = ((mul_34_17_n_5925 & mul_34_17_n_6101) | ((mul_34_17_n_5925 & mul_34_17_n_5924)
    | (mul_34_17_n_5924 & mul_34_17_n_6101)));
 assign mul_34_17_n_198 = (mul_34_17_n_6427 ^ mul_34_17_n_6100);
 assign mul_34_17_n_197 = (mul_34_17_n_6857 ^ mul_34_17_n_6075);
 assign mul_34_17_n_196 = (mul_34_17_n_6066 ^ mul_34_17_n_5327);
 assign mul_34_17_n_194 = ~mul_34_17_n_195;
 assign mul_34_17_n_195 = ((mul_34_17_n_5640 & mul_34_17_n_6063) | ((mul_34_17_n_5640 & mul_34_17_n_5972)
    | (mul_34_17_n_5972 & mul_34_17_n_6063)));
 assign mul_34_17_n_193 = (mul_34_17_n_6840 ^ mul_34_17_n_6041);
 assign mul_34_17_n_192 = (mul_34_17_n_6817 ^ mul_34_17_n_6037);
 assign mul_34_17_n_191 = (mul_34_17_n_6862 ^ mul_34_17_n_6035);
 assign mul_34_17_n_190 = (mul_34_17_n_5877 ^ mul_34_17_n_6025);
 assign mul_34_17_n_189 = (mul_34_17_n_6835 ^ mul_34_17_n_6020);
 assign mul_34_17_n_187 = ~mul_34_17_n_188;
 assign mul_34_17_n_188 = ((mul_34_17_n_6011 & mul_34_17_n_5763) | ((mul_34_17_n_6011 & mul_34_17_n_6018)
    | (mul_34_17_n_6018 & mul_34_17_n_5763)));
 assign mul_34_17_n_186 = (mul_34_17_n_7176 ^ mul_34_17_n_6003);
 assign mul_34_17_n_185 = (mul_34_17_n_6834 ^ mul_34_17_n_5977);
 assign mul_34_17_n_184 = (mul_34_17_n_6714 ^ mul_34_17_n_5973);
 assign mul_34_17_n_183 = (mul_34_17_n_6755 ^ mul_34_17_n_5957);
 assign mul_34_17_n_182 = (mul_34_17_n_6942 ^ mul_34_17_n_5947);
 assign mul_34_17_n_181 = (mul_34_17_n_6762 ^ mul_34_17_n_5926);
 assign mul_34_17_n_180 = (mul_34_17_n_6939 ^ mul_34_17_n_5802);
 assign mul_34_17_n_178 = ~mul_34_17_n_179;
 assign mul_34_17_n_179 = ((mul_34_17_n_5587 & mul_34_17_n_5781) | ((mul_34_17_n_5587 & mul_34_17_n_5572)
    | (mul_34_17_n_5572 & mul_34_17_n_5781)));
 assign mul_34_17_n_176 = ~mul_34_17_n_177;
 assign mul_34_17_n_177 = ((mul_34_17_n_5663 & mul_34_17_n_5759) | ((mul_34_17_n_5663 & mul_34_17_n_5664)
    | (mul_34_17_n_5664 & mul_34_17_n_5759)));
 assign mul_34_17_n_174 = ~mul_34_17_n_175;
 assign mul_34_17_n_175 = ((mul_34_17_n_5635 & mul_34_17_n_5747) | ((mul_34_17_n_5635 & mul_34_17_n_5508)
    | (mul_34_17_n_5508 & mul_34_17_n_5747)));
 assign mul_34_17_n_173 = (mul_34_17_n_6724 ^ mul_34_17_n_5741);
 assign mul_34_17_n_171 = ~mul_34_17_n_172;
 assign mul_34_17_n_172 = ((mul_34_17_n_5600 & mul_34_17_n_5735) | ((mul_34_17_n_5600 & mul_34_17_n_5546)
    | (mul_34_17_n_5546 & mul_34_17_n_5735)));
 assign mul_34_17_n_170 = (mul_34_17_n_6855 ^ mul_34_17_n_5725);
 assign mul_34_17_n_169 = (mul_34_17_n_6716 ^ mul_34_17_n_5715);
 assign mul_34_17_n_168 = (mul_34_17_n_6761 ^ mul_34_17_n_5713);
 assign mul_34_17_n_167 = (mul_34_17_n_6853 ^ mul_34_17_n_5683);
 assign mul_34_17_n_166 = (mul_34_17_n_6858 ^ mul_34_17_n_5672);
 assign mul_34_17_n_165 = (mul_34_17_n_6941 ^ mul_34_17_n_5654);
 assign mul_34_17_n_164 = (mul_34_17_n_7181 ^ mul_34_17_n_5645);
 assign mul_34_17_n_163 = (mul_34_17_n_6742 ^ mul_34_17_n_5644);
 assign mul_34_17_n_162 = (mul_34_17_n_6851 ^ mul_34_17_n_5638);
 assign mul_34_17_n_161 = (mul_34_17_n_6752 ^ mul_34_17_n_5623);
 assign mul_34_17_n_160 = (mul_34_17_n_6828 ^ mul_34_17_n_5607);
 assign mul_34_17_n_159 = (mul_34_17_n_6689 ^ mul_34_17_n_5556);
 assign mul_34_17_n_158 = (mul_34_17_n_6694 ^ mul_34_17_n_5550);
 assign mul_34_17_n_157 = (mul_34_17_n_6691 ^ mul_34_17_n_5547);
 assign mul_34_17_n_156 = (mul_34_17_n_6748 ^ mul_34_17_n_5524);
 assign mul_34_17_n_155 = (mul_34_17_n_6899 ^ mul_34_17_n_5504);
 assign mul_34_17_n_154 = (mul_34_17_n_5250 ^ mul_34_17_n_5448);
 assign mul_34_17_n_152 = (mul_34_17_n_5428 ^ mul_34_17_n_4886);
 assign mul_34_17_n_151 = (mul_34_17_n_6665 ^ mul_34_17_n_5425);
 assign mul_34_17_n_150 = (mul_34_17_n_5882 ^ mul_34_17_n_5415);
 assign mul_34_17_n_149 = (mul_34_17_n_5878 ^ mul_34_17_n_5414);
 assign mul_34_17_n_148 = (mul_34_17_n_5125 ^ mul_34_17_n_5881);
 assign mul_34_17_n_147 = (mul_34_17_n_5124 ^ mul_34_17_n_4845);
 assign mul_34_17_n_146 = (mul_34_17_n_5371 ^ mul_34_17_n_4815);
 assign mul_34_17_n_145 = (mul_34_17_n_5372 ^ mul_34_17_n_4811);
 assign mul_34_17_n_144 = (mul_34_17_n_5366 ^ mul_34_17_n_4804);
 assign mul_34_17_n_143 = (mul_34_17_n_5362 ^ mul_34_17_n_4801);
 assign mul_34_17_n_142 = (mul_34_17_n_5349 ^ mul_34_17_n_4778);
 assign mul_34_17_n_140 = ~mul_34_17_n_141;
 assign mul_34_17_n_141 = ((mul_34_17_n_4289 & mul_34_17_n_4769) | ((mul_34_17_n_4289 & mul_34_17_n_3427)
    | (mul_34_17_n_3427 & mul_34_17_n_4769)));
 assign mul_34_17_n_139 = (mul_34_17_n_4763 ^ mul_34_17_n_4107);
 assign mul_34_17_n_137 = ~mul_34_17_n_138;
 assign mul_34_17_n_138 = ((mul_34_17_n_4215 & mul_34_17_n_4762) | ((mul_34_17_n_4215 & mul_34_17_n_4223)
    | (mul_34_17_n_4223 & mul_34_17_n_4762)));
 assign mul_34_17_n_136 = (mul_34_17_n_5243 ^ mul_34_17_n_4758);
 assign mul_34_17_n_135 = (mul_34_17_n_5370 ^ mul_34_17_n_4728);
 assign mul_34_17_n_133 = ~mul_34_17_n_134;
 assign mul_34_17_n_134 = ((mul_34_17_n_4483 & mul_34_17_n_4715) | ((mul_34_17_n_4483 & mul_34_17_n_4486)
    | (mul_34_17_n_4486 & mul_34_17_n_4715)));
 assign mul_34_17_n_131 = ~mul_34_17_n_132;
 assign mul_34_17_n_132 = ((mul_34_17_n_4481 & mul_34_17_n_4712) | ((mul_34_17_n_4481 & mul_34_17_n_4159)
    | (mul_34_17_n_4159 & mul_34_17_n_4712)));
 assign mul_34_17_n_129 = ~mul_34_17_n_130;
 assign mul_34_17_n_130 = ((mul_34_17_n_4476 & mul_34_17_n_4710) | ((mul_34_17_n_4476 & mul_34_17_n_4123)
    | (mul_34_17_n_4123 & mul_34_17_n_4710)));
 assign mul_34_17_n_127 = ~mul_34_17_n_128;
 assign mul_34_17_n_128 = ((mul_34_17_n_3298 & mul_34_17_n_4695) | ((mul_34_17_n_3298 & mul_34_17_n_3301)
    | (mul_34_17_n_3301 & mul_34_17_n_4695)));
 assign mul_34_17_n_125 = ~mul_34_17_n_126;
 assign mul_34_17_n_126 = ((mul_34_17_n_4409 & mul_34_17_n_4693) | ((mul_34_17_n_4409 & mul_34_17_n_3365)
    | (mul_34_17_n_3365 & mul_34_17_n_4693)));
 assign mul_34_17_n_123 = ~mul_34_17_n_124;
 assign mul_34_17_n_124 = ((mul_34_17_n_4404 & mul_34_17_n_4691) | ((mul_34_17_n_4404 & mul_34_17_n_3610)
    | (mul_34_17_n_3610 & mul_34_17_n_4691)));
 assign mul_34_17_n_122 = (mul_34_17_n_5351 ^ mul_34_17_n_4684);
 assign mul_34_17_n_121 = (mul_34_17_n_5354 ^ mul_34_17_n_4682);
 assign mul_34_17_n_120 = (mul_34_17_n_5276 ^ mul_34_17_n_4671);
 assign mul_34_17_n_119 = (mul_34_17_n_5091 ^ mul_34_17_n_4667);
 assign mul_34_17_n_118 = (mul_34_17_n_5304 ^ mul_34_17_n_4660);
 assign mul_34_17_n_117 = (mul_34_17_n_5288 ^ mul_34_17_n_4656);
 assign mul_34_17_n_115 = (mul_34_17_n_5242 ^ mul_34_17_n_4637);
 assign mul_34_17_n_113 = ~mul_34_17_n_114;
 assign mul_34_17_n_114 = ((mul_34_17_n_4156 & mul_34_17_n_4623) | ((mul_34_17_n_4156 & mul_34_17_n_4157)
    | (mul_34_17_n_4157 & mul_34_17_n_4623)));
 assign mul_34_17_n_112 = (mul_34_17_n_5213 ^ mul_34_17_n_4614);
 assign mul_34_17_n_111 = (mul_34_17_n_5006 ^ mul_34_17_n_4613);
 assign mul_34_17_n_110 = (mul_34_17_n_4953 ^ mul_34_17_n_4609);
 assign mul_34_17_n_108 = ~mul_34_17_n_109;
 assign mul_34_17_n_109 = ((mul_34_17_n_4278 & mul_34_17_n_4608) | ((mul_34_17_n_4278 & mul_34_17_n_4280)
    | (mul_34_17_n_4280 & mul_34_17_n_4608)));
 assign mul_34_17_n_107 = (mul_34_17_n_5227 ^ mul_34_17_n_4601);
 assign mul_34_17_n_105 = ~mul_34_17_n_106;
 assign mul_34_17_n_106 = ((mul_34_17_n_3601 & mul_34_17_n_4594) | ((mul_34_17_n_3601 & mul_34_17_n_3625)
    | (mul_34_17_n_3625 & mul_34_17_n_4594)));
 assign mul_34_17_n_103 = ~mul_34_17_n_104;
 assign mul_34_17_n_104 = ((mul_34_17_n_4399 & mul_34_17_n_4588) | ((mul_34_17_n_4399 & mul_34_17_n_4036)
    | (mul_34_17_n_4036 & mul_34_17_n_4588)));
 assign mul_34_17_n_102 = (mul_34_17_n_4916 ^ mul_34_17_n_4586);
 assign mul_34_17_n_101 = (mul_34_17_n_5214 ^ mul_34_17_n_4585);
 assign mul_34_17_n_99 = ~mul_34_17_n_100;
 assign mul_34_17_n_100 = ((mul_34_17_n_3261 & mul_34_17_n_4571) | ((mul_34_17_n_3261 & mul_34_17_n_3651)
    | (mul_34_17_n_3651 & mul_34_17_n_4571)));
 assign mul_34_17_n_98 = (mul_34_17_n_5027 ^ mul_34_17_n_4548);
 assign mul_34_17_n_97 = (mul_34_17_n_5041 ^ mul_34_17_n_4541);
 assign mul_34_17_n_96 = (mul_34_17_n_4928 ^ mul_34_17_n_4410);
 assign mul_34_17_n_95 = (mul_34_17_n_5384 ^ mul_34_17_n_4371);
 assign mul_34_17_n_94 = (mul_34_17_n_5266 ^ mul_34_17_n_4323);
 assign mul_34_17_n_93 = (mul_34_17_n_5310 ^ mul_34_17_n_4302);
 assign mul_34_17_n_92 = (mul_34_17_n_5008 ^ mul_34_17_n_4268);
 assign mul_34_17_n_91 = (mul_34_17_n_5323 ^ mul_34_17_n_4226);
 assign mul_34_17_n_89 = ~mul_34_17_n_90;
 assign mul_34_17_n_90 = ((mul_34_17_n_3385 & mul_34_17_n_3733) | ((mul_34_17_n_3385 & mul_34_17_n_4211)
    | (mul_34_17_n_4211 & mul_34_17_n_3733)));
 assign mul_34_17_n_88 = (mul_34_17_n_5012 ^ mul_34_17_n_4207);
 assign mul_34_17_n_87 = (mul_34_17_n_5286 ^ mul_34_17_n_4174);
 assign mul_34_17_n_85 = ~mul_34_17_n_86;
 assign mul_34_17_n_86 = ((mul_34_17_n_3624 & mul_34_17_n_3759) | ((mul_34_17_n_3624 & mul_34_17_n_4142)
    | (mul_34_17_n_4142 & mul_34_17_n_3759)));
 assign mul_34_17_n_84 = (mul_34_17_n_5212 ^ mul_34_17_n_4125);
 assign mul_34_17_n_83 = (mul_34_17_n_5211 ^ mul_34_17_n_4121);
 assign mul_34_17_n_82 = (mul_34_17_n_5334 ^ mul_34_17_n_4104);
 assign mul_34_17_n_81 = (mul_34_17_n_5317 ^ mul_34_17_n_4082);
 assign mul_34_17_n_80 = (mul_34_17_n_5350 ^ mul_34_17_n_4073);
 assign mul_34_17_n_79 = (mul_34_17_n_5016 ^ mul_34_17_n_4051);
 assign mul_34_17_n_77 = ~mul_34_17_n_78;
 assign mul_34_17_n_78 = ~(mul_34_17_n_4049 | mul_34_17_n_3967);
 assign mul_34_17_n_75 = ~mul_34_17_n_76;
 assign mul_34_17_n_76 = ((mul_34_17_n_4037 & mul_34_17_n_3723) | ((mul_34_17_n_4037 & mul_34_17_n_3582)
    | (mul_34_17_n_3582 & mul_34_17_n_3723)));
 assign mul_34_17_n_73 = ~mul_34_17_n_74;
 assign mul_34_17_n_74 = ((mul_34_17_n_4030 & mul_34_17_n_3817) | ((mul_34_17_n_4030 & mul_34_17_n_4029)
    | (mul_34_17_n_4029 & mul_34_17_n_3817)));
 assign mul_34_17_n_72 = (mul_34_17_n_5430 ^ mul_34_17_n_3980);
 assign mul_34_17_n_71 = (mul_34_17_n_5435 ^ mul_34_17_n_3977);
 assign mul_34_17_n_69 = ~mul_34_17_n_70;
 assign mul_34_17_n_70 = ((mul_34_17_n_3158 & mul_34_17_n_3976) | ((mul_34_17_n_3158 & mul_34_17_n_3256)
    | (mul_34_17_n_3256 & mul_34_17_n_3976)));
 assign mul_34_17_n_67 = ~mul_34_17_n_68;
 assign mul_34_17_n_68 = ~(mul_34_17_n_3975 & mul_34_17_n_3932);
 assign mul_34_17_n_66 = (mul_34_17_n_5315 ^ mul_34_17_n_3925);
 assign mul_34_17_n_65 = (mul_34_17_n_5271 ^ mul_34_17_n_3924);
 assign mul_34_17_n_64 = (mul_34_17_n_5291 ^ mul_34_17_n_3919);
 assign mul_34_17_n_63 = (mul_34_17_n_5249 ^ mul_34_17_n_3915);
 assign mul_34_17_n_62 = (mul_34_17_n_5382 ^ mul_34_17_n_3912);
 assign mul_34_17_n_61 = (mul_34_17_n_5045 ^ mul_34_17_n_3909);
 assign mul_34_17_n_59 = ~mul_34_17_n_60;
 assign mul_34_17_n_60 = ((mul_34_17_n_3058 & mul_34_17_n_3899) | ((mul_34_17_n_3058 & mul_34_17_n_3575)
    | (mul_34_17_n_3575 & mul_34_17_n_3899)));
 assign mul_34_17_n_58 = (mul_34_17_n_5270 ^ mul_34_17_n_3887);
 assign mul_34_17_n_56 = ~mul_34_17_n_57;
 assign mul_34_17_n_57 = ((mul_34_17_n_3251 & mul_34_17_n_3880) | ((mul_34_17_n_3251 & mul_34_17_n_3156)
    | (mul_34_17_n_3156 & mul_34_17_n_3880)));
 assign mul_34_17_n_55 = (mul_34_17_n_5023 ^ mul_34_17_n_3873);
 assign mul_34_17_n_54 = (mul_34_17_n_5033 ^ mul_34_17_n_3864);
 assign mul_34_17_n_53 = (mul_34_17_n_5373 ^ mul_34_17_n_3835);
 assign mul_34_17_n_52 = (mul_34_17_n_5009 ^ mul_34_17_n_3832);
 assign mul_34_17_n_51 = (mul_34_17_n_5230 ^ mul_34_17_n_3818);
 assign mul_34_17_n_49 = ~mul_34_17_n_50;
 assign mul_34_17_n_50 = ((mul_34_17_n_3440 & mul_34_17_n_3813) | ((mul_34_17_n_3440 & mul_34_17_n_3343)
    | (mul_34_17_n_3343 & mul_34_17_n_3813)));
 assign mul_34_17_n_48 = (mul_34_17_n_5328 ^ mul_34_17_n_3810);
 assign mul_34_17_n_46 = ~mul_34_17_n_47;
 assign mul_34_17_n_47 = ((mul_34_17_n_3485 & mul_34_17_n_3800) | ((mul_34_17_n_3485 & mul_34_17_n_3487)
    | (mul_34_17_n_3487 & mul_34_17_n_3800)));
 assign mul_34_17_n_45 = (mul_34_17_n_5256 ^ mul_34_17_n_3791);
 assign mul_34_17_n_43 = ~mul_34_17_n_44;
 assign mul_34_17_n_44 = ((mul_34_17_n_3448 & mul_34_17_n_3787) | ((mul_34_17_n_3448 & mul_34_17_n_3449)
    | (mul_34_17_n_3449 & mul_34_17_n_3787)));
 assign mul_34_17_n_42 = (mul_34_17_n_5225 ^ mul_34_17_n_3785);
 assign mul_34_17_n_41 = (mul_34_17_n_5289 ^ mul_34_17_n_3782);
 assign mul_34_17_n_40 = (mul_34_17_n_5074 ^ mul_34_17_n_3754);
 assign mul_34_17_n_39 = (mul_34_17_n_5073 ^ mul_34_17_n_3729);
 assign mul_34_17_n_38 = (mul_34_17_n_5287 ^ mul_34_17_n_3725);
 assign mul_34_17_n_37 = (mul_34_17_n_5071 ^ mul_34_17_n_3717);
 assign mul_34_17_n_36 = (mul_34_17_n_4920 ^ mul_34_17_n_3714);
 assign mul_34_17_n_35 = (mul_34_17_n_4952 ^ mul_34_17_n_3713);
 assign mul_34_17_n_34 = (mul_34_17_n_4924 ^ mul_34_17_n_3692);
 assign mul_34_17_n_32 = ~mul_34_17_n_33;
 assign mul_34_17_n_33 = ((mul_34_17_n_3430 & mul_34_17_n_3677) | ((mul_34_17_n_3430 & mul_34_17_n_3432)
    | (mul_34_17_n_3432 & mul_34_17_n_3677)));
 assign mul_34_17_n_31 = (mul_34_17_n_5010 ^ mul_34_17_n_3675);
 assign mul_34_17_n_30 = (mul_34_17_n_5036 ^ mul_34_17_n_3673);
 assign mul_34_17_n_29 = (mul_34_17_n_5079 ^ mul_34_17_n_3667);
 assign mul_34_17_n_28 = (mul_34_17_n_5378 ^ mul_34_17_n_3598);
 assign mul_34_17_n_27 = (mul_34_17_n_5014 ^ mul_34_17_n_3571);
 assign mul_34_17_n_26 = (mul_34_17_n_5068 ^ mul_34_17_n_3562);
 assign mul_34_17_n_25 = (mul_34_17_n_5001 ^ mul_34_17_n_3546);
 assign mul_34_17_n_24 = (mul_34_17_n_5231 ^ mul_34_17_n_3530);
 assign mul_34_17_n_23 = (mul_34_17_n_4987 ^ mul_34_17_n_3499);
 assign mul_34_17_n_22 = (mul_34_17_n_4943 ^ mul_34_17_n_3482);
 assign mul_34_17_n_21 = (mul_34_17_n_4963 ^ mul_34_17_n_3478);
 assign mul_34_17_n_20 = (mul_34_17_n_5002 ^ mul_34_17_n_3473);
 assign mul_34_17_n_19 = (mul_34_17_n_4932 ^ mul_34_17_n_3471);
 assign mul_34_17_n_18 = (mul_34_17_n_4964 ^ mul_34_17_n_3367);
 assign mul_34_17_n_17 = (mul_34_17_n_5087 ^ mul_34_17_n_3362);
 assign mul_34_17_n_16 = (mul_34_17_n_5238 ^ mul_34_17_n_3353);
 assign mul_34_17_n_15 = (mul_34_17_n_5240 ^ mul_34_17_n_3306);
 assign mul_34_17_n_14 = (mul_34_17_n_5255 ^ mul_34_17_n_3254);
 assign mul_34_17_n_13 = (mul_34_17_n_4930 ^ mul_34_17_n_3209);
 assign mul_34_17_n_12 = (mul_34_17_n_5092 ^ mul_34_17_n_3193);
 assign mul_34_17_n_11 = (mul_34_17_n_4925 ^ mul_34_17_n_3188);
 assign mul_34_17_n_10 = (mul_34_17_n_4922 ^ mul_34_17_n_3184);
 assign mul_34_17_n_8 = ~mul_34_17_n_9;
 assign mul_34_17_n_9 = ((mul_34_17_n_3182 & mul_34_17_n_3173) | ((mul_34_17_n_3182 & mul_34_17_n_3174)
    | (mul_34_17_n_3174 & mul_34_17_n_3173)));
 assign mul_34_17_n_7 = (mul_34_17_n_5314 ^ mul_34_17_n_3150);
 assign mul_34_17_n_6 = (mul_34_17_n_5126 ^ mul_34_17_n_3059);
 assign mul_34_17_n_5 = (mul_34_17_n_2860 ^ mul_34_17_n_2949);
 assign mul_34_17_n_4 = (mul_34_17_n_2850 ^ mul_34_17_n_2938);
 assign mul_34_17_n_3 = (mul_34_17_n_4913 ^ mul_34_17_n_2838);
 assign mul_34_17_n_2 = (mul_34_17_n_5296 ^ mul_34_17_n_2823);
 assign mul_34_17_n_1 = (mul_34_17_n_4933 ^ mul_34_17_n_2816);
 assign mul_34_17_n_0 = (mul_34_17_n_8822 ^ mul_34_17_n_225);
 assign mul_34_17_n_11272 = ~(mul_34_17_n_9716 ^ (mul_34_17_n_9528 ^ (mul_34_17_n_9280 ^ mul_34_17_n_9717)));
 assign mul_34_17_n_11274 = (mul_34_17_n_9487 ^ mul_34_17_n_11273);
 assign mul_34_17_n_11273 = (mul_34_17_n_9464 ^ mul_34_17_n_9265);
 assign mul_34_17_n_11276 = (mul_34_17_n_9485 ^ mul_34_17_n_11275);
 assign mul_34_17_n_11275 = (mul_34_17_n_9470 ^ mul_34_17_n_9334);
 assign mul_34_17_n_11278 = (mul_34_17_n_9332 ^ mul_34_17_n_11277);
 assign mul_34_17_n_11277 = ~(mul_34_17_n_9466 ^ mul_34_17_n_9160);
 assign mul_34_17_n_11280 = (mul_34_17_n_355 ^ mul_34_17_n_11279);
 assign mul_34_17_n_11279 = (mul_34_17_n_9094 ^ mul_34_17_n_9100);
 assign mul_34_17_n_11282 = (mul_34_17_n_9172 ^ mul_34_17_n_11281);
 assign mul_34_17_n_11281 = ~(mul_34_17_n_278 ^ mul_34_17_n_9166);
 assign mul_34_17_n_11284 = (mul_34_17_n_276 ^ mul_34_17_n_11283);
 assign mul_34_17_n_11283 = ~(mul_34_17_n_9354 ^ mul_34_17_n_9352);
 assign mul_34_17_n_11286 = (mul_34_17_n_286 ^ mul_34_17_n_11285);
 assign mul_34_17_n_11285 = (mul_34_17_n_11320 ^ mul_34_17_n_9158);
 assign mul_34_17_n_11288 = (mul_34_17_n_9493 ^ mul_34_17_n_11287);
 assign mul_34_17_n_11287 = (mul_34_17_n_9356 ^ mul_34_17_n_11316);
 assign mul_34_17_n_11290 = ~mul_34_17_n_11289;
 assign mul_34_17_n_11289 = ((mul_34_17_n_9483 & mul_34_17_n_9196) | ((mul_34_17_n_9483 & mul_34_17_n_9333)
    | (mul_34_17_n_9333 & mul_34_17_n_9196)));
 assign mul_34_17_n_11292 = ((mul_34_17_n_9271 & mul_34_17_n_11291) | ((mul_34_17_n_9271 & mul_34_17_n_8992)
    | (mul_34_17_n_8992 & mul_34_17_n_11291)));
 assign mul_34_17_n_11291 = ~(mul_34_17_n_9006 ^ mul_34_17_n_8492);
 assign mul_34_17_n_11294 = ~mul_34_17_n_11293;
 assign mul_34_17_n_11293 = ((mul_34_17_n_9268 & mul_34_17_n_264) | ((mul_34_17_n_9268 & mul_34_17_n_9260)
    | (mul_34_17_n_9260 & mul_34_17_n_264)));
 assign mul_34_17_n_11296 = ~mul_34_17_n_11295;
 assign mul_34_17_n_11295 = ((mul_34_17_n_285 & mul_34_17_n_9191) | ((mul_34_17_n_285 & mul_34_17_n_9190)
    | (mul_34_17_n_9190 & mul_34_17_n_9191)));
 assign mul_34_17_n_11298 = (mul_34_17_n_9200 ^ mul_34_17_n_11297);
 assign mul_34_17_n_11297 = (mul_34_17_n_11346 ^ mul_34_17_n_9104);
 assign mul_34_17_n_11300 = (mul_34_17_n_9031 ^ mul_34_17_n_11299);
 assign mul_34_17_n_11299 = (mul_34_17_n_8993 ^ mul_34_17_n_9017);
 assign mul_34_17_n_11302 = ((mul_34_17_n_9005 & mul_34_17_n_11301) | ((mul_34_17_n_9005 & mul_34_17_n_8851)
    | (mul_34_17_n_8851 & mul_34_17_n_11301)));
 assign mul_34_17_n_11301 = (mul_34_17_n_8850 ^ mul_34_17_n_8598);
 assign mul_34_17_n_11304 = (mul_34_17_n_268 ^ mul_34_17_n_11303);
 assign mul_34_17_n_11303 = (mul_34_17_n_9089 ^ mul_34_17_n_8984);
 assign mul_34_17_n_11306 = (mul_34_17_n_274 ^ mul_34_17_n_11305);
 assign mul_34_17_n_11305 = ~(mul_34_17_n_8838 ^ mul_34_17_n_9014);
 assign mul_34_17_n_11308 = ~mul_34_17_n_11307;
 assign mul_34_17_n_11307 = ((mul_34_17_n_362 & mul_34_17_n_9277) | ((mul_34_17_n_362 & mul_34_17_n_8732)
    | (mul_34_17_n_8732 & mul_34_17_n_9277)));
 assign mul_34_17_n_11310 = (mul_34_17_n_9007 ^ mul_34_17_n_11309);
 assign mul_34_17_n_11309 = (mul_34_17_n_11348 ^ mul_34_17_n_8730);
 assign mul_34_17_n_11312 = (mul_34_17_n_273 ^ mul_34_17_n_11311);
 assign mul_34_17_n_11311 = ~(mul_34_17_n_8834 ^ mul_34_17_n_8724);
 assign mul_34_17_n_11314 = (mul_34_17_n_8938 ^ mul_34_17_n_11313);
 assign mul_34_17_n_11313 = (mul_34_17_n_8744 ^ mul_34_17_n_8537);
 assign mul_34_17_n_11316 = (mul_34_17_n_8682 ^ mul_34_17_n_11315);
 assign mul_34_17_n_11315 = (mul_34_17_n_8664 ^ mul_34_17_n_8346);
 assign mul_34_17_n_11318 = (mul_34_17_n_8773 ^ mul_34_17_n_11317);
 assign mul_34_17_n_11317 = ~(mul_34_17_n_8739 ^ mul_34_17_n_8140);
 assign mul_34_17_n_11320 = (mul_34_17_n_8782 ^ mul_34_17_n_11319);
 assign mul_34_17_n_11319 = ~(mul_34_17_n_8766 ^ mul_34_17_n_8252);
 assign mul_34_17_n_11322 = (mul_34_17_n_8922 ^ mul_34_17_n_11321);
 assign mul_34_17_n_11321 = ~(mul_34_17_n_8609 ^ mul_34_17_n_8723);
 assign mul_34_17_n_11324 = (mul_34_17_n_8777 ^ mul_34_17_n_11323);
 assign mul_34_17_n_11323 = (mul_34_17_n_8525 ^ mul_34_17_n_11378);
 assign mul_34_17_n_11326 = (mul_34_17_n_8524 ^ mul_34_17_n_11325);
 assign mul_34_17_n_11325 = ~(mul_34_17_n_8227 ^ mul_34_17_n_8485);
 assign mul_34_17_n_11328 = ((mul_34_17_n_11394 & mul_34_17_n_11327) | ((mul_34_17_n_11394 & mul_34_17_n_8036)
    | (mul_34_17_n_8036 & mul_34_17_n_11327)));
 assign mul_34_17_n_11327 = (mul_34_17_n_8132 ^ mul_34_17_n_7437);
 assign mul_34_17_n_11330 = (mul_34_17_n_224 ^ mul_34_17_n_11329);
 assign mul_34_17_n_11329 = ~(mul_34_17_n_11481 ^ mul_34_17_n_8224);
 assign mul_34_17_n_11332 = (mul_34_17_n_233 ^ mul_34_17_n_11331);
 assign mul_34_17_n_11331 = ~(mul_34_17_n_7998 ^ mul_34_17_n_8253);
 assign mul_34_17_n_11334 = (mul_34_17_n_8153 ^ mul_34_17_n_11333);
 assign mul_34_17_n_11333 = ~(mul_34_17_n_8007 ^ mul_34_17_n_8028);
 assign mul_34_17_n_11336 = (mul_34_17_n_159 ^ mul_34_17_n_11335);
 assign mul_34_17_n_11335 = (mul_34_17_n_11472 ^ mul_34_17_n_11476);
 assign mul_34_17_n_11338 = (mul_34_17_n_8003 ^ mul_34_17_n_11337);
 assign mul_34_17_n_11337 = (mul_34_17_n_11629 ^ mul_34_17_n_182);
 assign mul_34_17_n_11340 = (mul_34_17_n_8019 ^ mul_34_17_n_11339);
 assign mul_34_17_n_11339 = (mul_34_17_n_11404 ^ mul_34_17_n_11414);
 assign mul_34_17_n_11342 = (mul_34_17_n_7492 ^ mul_34_17_n_11341);
 assign mul_34_17_n_11341 = (mul_34_17_n_11466 ^ mul_34_17_n_7986);
 assign mul_34_17_n_11344 = (mul_34_17_n_7900 ^ mul_34_17_n_11343);
 assign mul_34_17_n_11343 = (mul_34_17_n_11406 ^ mul_34_17_n_11479);
 assign mul_34_17_n_11346 = (mul_34_17_n_7483 ^ mul_34_17_n_11345);
 assign mul_34_17_n_11345 = ~(mul_34_17_n_7853 ^ mul_34_17_n_7832);
 assign mul_34_17_n_11348 = (mul_34_17_n_7700 ^ mul_34_17_n_11347);
 assign mul_34_17_n_11347 = ~(mul_34_17_n_11474 ^ mul_34_17_n_11468);
 assign mul_34_17_n_11350 = (mul_34_17_n_7146 ^ mul_34_17_n_11349);
 assign mul_34_17_n_11349 = ~(mul_34_17_n_7500 ^ mul_34_17_n_6896);
 assign mul_34_17_n_11352 = (mul_34_17_n_7932 ^ mul_34_17_n_11351);
 assign mul_34_17_n_11351 = ~(mul_34_17_n_7545 ^ mul_34_17_n_7544);
 assign mul_34_17_n_11354 = (mul_34_17_n_7579 ^ mul_34_17_n_11353);
 assign mul_34_17_n_11353 = ~(mul_34_17_n_7503 ^ mul_34_17_n_7501);
 assign mul_34_17_n_11356 = (mul_34_17_n_7517 ^ mul_34_17_n_11355);
 assign mul_34_17_n_11355 = (mul_34_17_n_7413 ^ mul_34_17_n_7682);
 assign mul_34_17_n_11358 = (mul_34_17_n_7534 ^ mul_34_17_n_11357);
 assign mul_34_17_n_11357 = ~(mul_34_17_n_7679 ^ mul_34_17_n_7408);
 assign mul_34_17_n_11360 = (mul_34_17_n_7537 ^ mul_34_17_n_11359);
 assign mul_34_17_n_11359 = ~(mul_34_17_n_7431 ^ mul_34_17_n_7407);
 assign mul_34_17_n_11362 = (mul_34_17_n_7779 ^ mul_34_17_n_11361);
 assign mul_34_17_n_11361 = (mul_34_17_n_7724 ^ mul_34_17_n_7511);
 assign mul_34_17_n_11364 = (mul_34_17_n_7533 ^ mul_34_17_n_11363);
 assign mul_34_17_n_11363 = ~(mul_34_17_n_7433 ^ mul_34_17_n_7418);
 assign mul_34_17_n_11366 = (mul_34_17_n_173 ^ mul_34_17_n_11365);
 assign mul_34_17_n_11365 = ~(mul_34_17_n_7438 ^ mul_34_17_n_7420);
 assign mul_34_17_n_11368 = (mul_34_17_n_7469 ^ mul_34_17_n_11367);
 assign mul_34_17_n_11367 = ~(mul_34_17_n_7440 ^ mul_34_17_n_7425);
 assign mul_34_17_n_11370 = (mul_34_17_n_6798 ^ mul_34_17_n_11369);
 assign mul_34_17_n_11369 = ~(mul_34_17_n_7075 ^ mul_34_17_n_6340);
 assign mul_34_17_n_11372 = (mul_34_17_n_6789 ^ mul_34_17_n_11371);
 assign mul_34_17_n_11371 = ~(mul_34_17_n_7291 ^ mul_34_17_n_6497);
 assign mul_34_17_n_11374 = (mul_34_17_n_7542 ^ mul_34_17_n_11373);
 assign mul_34_17_n_11373 = ~(mul_34_17_n_7058 ^ mul_34_17_n_6454);
 assign mul_34_17_n_11376 = (mul_34_17_n_7473 ^ mul_34_17_n_11375);
 assign mul_34_17_n_11375 = ~(mul_34_17_n_7057 ^ mul_34_17_n_7050);
 assign mul_34_17_n_11378 = (mul_34_17_n_7711 ^ mul_34_17_n_11377);
 assign mul_34_17_n_11377 = ~(mul_34_17_n_7292 ^ mul_34_17_n_6893);
 assign mul_34_17_n_11380 = (mul_34_17_n_7491 ^ mul_34_17_n_11379);
 assign mul_34_17_n_11379 = ~(mul_34_17_n_7051 ^ mul_34_17_n_7056);
 assign mul_34_17_n_11382 = (mul_34_17_n_6655 ^ mul_34_17_n_11381);
 assign mul_34_17_n_11381 = (mul_34_17_n_6581 ^ mul_34_17_n_6584);
 assign mul_34_17_n_11384 = (mul_34_17_n_6382 ^ mul_34_17_n_11383);
 assign mul_34_17_n_11383 = (mul_34_17_n_6273 ^ mul_34_17_n_6271);
 assign mul_34_17_n_11386 = (mul_34_17_n_6358 ^ mul_34_17_n_11385);
 assign mul_34_17_n_11385 = ~(mul_34_17_n_6320 ^ mul_34_17_n_6322);
 assign mul_34_17_n_11388 = (mul_34_17_n_66 ^ mul_34_17_n_11387);
 assign mul_34_17_n_11387 = (mul_34_17_n_117 ^ mul_34_17_n_65);
 assign mul_34_17_n_11390 = (mul_34_17_n_6365 ^ mul_34_17_n_11389);
 assign mul_34_17_n_11389 = (mul_34_17_n_6325 ^ mul_34_17_n_6319);
 assign mul_34_17_n_11392 = (mul_34_17_n_6637 ^ mul_34_17_n_11391);
 assign mul_34_17_n_11391 = (mul_34_17_n_41 ^ mul_34_17_n_38);
 assign mul_34_17_n_11394 = (mul_34_17_n_12 ^ mul_34_17_n_11393);
 assign mul_34_17_n_11393 = ~(mul_34_17_n_17 ^ mul_34_17_n_5122);
 assign mul_34_17_n_11396 = (mul_34_17_n_23 ^ mul_34_17_n_11395);
 assign mul_34_17_n_11395 = (mul_34_17_n_6275 ^ mul_34_17_n_18);
 assign mul_34_17_n_11398 = (mul_34_17_n_101 ^ mul_34_17_n_11397);
 assign mul_34_17_n_11397 = (mul_34_17_n_111 ^ mul_34_17_n_112);
 assign mul_34_17_n_11400 = (mul_34_17_n_6650 ^ mul_34_17_n_11399);
 assign mul_34_17_n_11399 = ~(mul_34_17_n_6560 ^ mul_34_17_n_5133);
 assign mul_34_17_n_11402 = (mul_34_17_n_6657 ^ mul_34_17_n_11401);
 assign mul_34_17_n_11401 = ~(mul_34_17_n_6019 ^ mul_34_17_n_6613);
 assign mul_34_17_n_11404 = (mul_34_17_n_6671 ^ mul_34_17_n_11403);
 assign mul_34_17_n_11403 = (mul_34_17_n_6550 ^ mul_34_17_n_6548);
 assign mul_34_17_n_11406 = (mul_34_17_n_6381 ^ mul_34_17_n_11405);
 assign mul_34_17_n_11405 = ~(mul_34_17_n_6281 ^ mul_34_17_n_6280);
 assign mul_34_17_n_11408 = (mul_34_17_n_6374 ^ mul_34_17_n_11407);
 assign mul_34_17_n_11407 = ~(mul_34_17_n_6289 ^ mul_34_17_n_6287);
 assign mul_34_17_n_11410 = (mul_34_17_n_6640 ^ mul_34_17_n_11409);
 assign mul_34_17_n_11409 = ~(mul_34_17_n_6533 ^ mul_34_17_n_6534);
 assign mul_34_17_n_11412 = (mul_34_17_n_6371 ^ mul_34_17_n_11411);
 assign mul_34_17_n_11411 = (mul_34_17_n_6291 ^ mul_34_17_n_6294);
 assign mul_34_17_n_11414 = (mul_34_17_n_6668 ^ mul_34_17_n_11413);
 assign mul_34_17_n_11413 = (mul_34_17_n_6557 ^ mul_34_17_n_6556);
 assign mul_34_17_n_11416 = (mul_34_17_n_154 ^ mul_34_17_n_11415);
 assign mul_34_17_n_11415 = ~(mul_34_17_n_6571 ^ mul_34_17_n_6570);
 assign mul_34_17_n_11418 = (mul_34_17_n_6632 ^ mul_34_17_n_11417);
 assign mul_34_17_n_11417 = ~(mul_34_17_n_6536 ^ mul_34_17_n_6539);
 assign mul_34_17_n_11420 = (mul_34_17_n_6232 ^ mul_34_17_n_11419);
 assign mul_34_17_n_11419 = (mul_34_17_n_13 ^ mul_34_17_n_96);
 assign mul_34_17_n_11422 = (mul_34_17_n_6300 ^ mul_34_17_n_11421);
 assign mul_34_17_n_11421 = (mul_34_17_n_63 ^ mul_34_17_n_118);
 assign mul_34_17_n_11424 = (mul_34_17_n_6245 ^ mul_34_17_n_11423);
 assign mul_34_17_n_11423 = ~(mul_34_17_n_6210 ^ mul_34_17_n_6154);
 assign mul_34_17_n_11426 = (mul_34_17_n_6588 ^ mul_34_17_n_11425);
 assign mul_34_17_n_11425 = ~(mul_34_17_n_6507 ^ mul_34_17_n_6484);
 assign mul_34_17_n_11428 = (mul_34_17_n_6530 ^ mul_34_17_n_11427);
 assign mul_34_17_n_11427 = (mul_34_17_n_6452 ^ mul_34_17_n_6500);
 assign mul_34_17_n_11430 = (mul_34_17_n_6282 ^ mul_34_17_n_11429);
 assign mul_34_17_n_11429 = ~(mul_34_17_n_79 ^ mul_34_17_n_97);
 assign mul_34_17_n_11432 = (mul_34_17_n_6617 ^ mul_34_17_n_11431);
 assign mul_34_17_n_11431 = ~(mul_34_17_n_6505 ^ mul_34_17_n_6480);
 assign mul_34_17_n_11434 = (mul_34_17_n_6800 ^ mul_34_17_n_11433);
 assign mul_34_17_n_11433 = (mul_34_17_n_6156 ^ mul_34_17_n_6174);
 assign mul_34_17_n_11436 = (mul_34_17_n_6385 ^ mul_34_17_n_11435);
 assign mul_34_17_n_11435 = (mul_34_17_n_6254 ^ mul_34_17_n_6259);
 assign mul_34_17_n_11438 = (mul_34_17_n_5141 ^ mul_34_17_n_11437);
 assign mul_34_17_n_11437 = (mul_34_17_n_25 ^ mul_34_17_n_6237);
 assign mul_34_17_n_11440 = (mul_34_17_n_6559 ^ mul_34_17_n_11439);
 assign mul_34_17_n_11439 = ~(mul_34_17_n_6458 ^ mul_34_17_n_6498);
 assign mul_34_17_n_11442 = (mul_34_17_n_6563 ^ mul_34_17_n_11441);
 assign mul_34_17_n_11441 = ~(mul_34_17_n_6503 ^ mul_34_17_n_6459);
 assign mul_34_17_n_11444 = (mul_34_17_n_6396 ^ mul_34_17_n_11443);
 assign mul_34_17_n_11443 = ~(mul_34_17_n_88 ^ mul_34_17_n_98);
 assign mul_34_17_n_11446 = (mul_34_17_n_6256 ^ mul_34_17_n_11445);
 assign mul_34_17_n_11445 = (mul_34_17_n_6206 ^ mul_34_17_n_6181);
 assign mul_34_17_n_11448 = (mul_34_17_n_6221 ^ mul_34_17_n_11447);
 assign mul_34_17_n_11447 = (mul_34_17_n_6191 ^ mul_34_17_n_6214);
 assign mul_34_17_n_11450 = (mul_34_17_n_6366 ^ mul_34_17_n_11449);
 assign mul_34_17_n_11449 = ~(mul_34_17_n_6306 ^ mul_34_17_n_6313);
 assign mul_34_17_n_11452 = (mul_34_17_n_6380 ^ mul_34_17_n_11451);
 assign mul_34_17_n_11451 = ~(mul_34_17_n_6284 ^ mul_34_17_n_6285);
 assign mul_34_17_n_11454 = (mul_34_17_n_7148 ^ mul_34_17_n_11453);
 assign mul_34_17_n_11453 = ~(mul_34_17_n_5708 ^ mul_34_17_n_7);
 assign mul_34_17_n_11456 = (mul_34_17_n_42 ^ mul_34_17_n_11455);
 assign mul_34_17_n_11455 = ~(mul_34_17_n_48 ^ mul_34_17_n_24);
 assign mul_34_17_n_11458 = (mul_34_17_n_6620 ^ mul_34_17_n_11457);
 assign mul_34_17_n_11457 = ~(mul_34_17_n_6478 ^ mul_34_17_n_6510);
 assign mul_34_17_n_11460 = (mul_34_17_n_6315 ^ mul_34_17_n_11459);
 assign mul_34_17_n_11459 = (mul_34_17_n_6479 ^ mul_34_17_n_6518);
 assign mul_34_17_n_11462 = (mul_34_17_n_6332 ^ mul_34_17_n_11461);
 assign mul_34_17_n_11461 = (mul_34_17_n_6192 ^ mul_34_17_n_6153);
 assign mul_34_17_n_11464 = (mul_34_17_n_6619 ^ mul_34_17_n_11463);
 assign mul_34_17_n_11463 = ~(mul_34_17_n_6526 ^ mul_34_17_n_6472);
 assign mul_34_17_n_11466 = (mul_34_17_n_6628 ^ mul_34_17_n_11465);
 assign mul_34_17_n_11465 = ~(mul_34_17_n_6160 ^ mul_34_17_n_6163);
 assign mul_34_17_n_11468 = (mul_34_17_n_6608 ^ mul_34_17_n_11467);
 assign mul_34_17_n_11467 = ~(mul_34_17_n_6513 ^ mul_34_17_n_6469);
 assign mul_34_17_n_11470 = (mul_34_17_n_142 ^ mul_34_17_n_11469);
 assign mul_34_17_n_11469 = (mul_34_17_n_34 ^ mul_34_17_n_122);
 assign mul_34_17_n_11472 = (mul_34_17_n_6266 ^ mul_34_17_n_11471);
 assign mul_34_17_n_11471 = (mul_34_17_n_6189 ^ mul_34_17_n_6205);
 assign mul_34_17_n_11474 = (mul_34_17_n_6606 ^ mul_34_17_n_11473);
 assign mul_34_17_n_11473 = ~(mul_34_17_n_6522 ^ mul_34_17_n_6467);
 assign mul_34_17_n_11476 = (mul_34_17_n_6267 ^ mul_34_17_n_11475);
 assign mul_34_17_n_11475 = (mul_34_17_n_6204 ^ mul_34_17_n_6164);
 assign mul_34_17_n_11478 = (mul_34_17_n_6623 ^ mul_34_17_n_11477);
 assign mul_34_17_n_11477 = ~(mul_34_17_n_6514 ^ mul_34_17_n_6474);
 assign mul_34_17_n_11479 = (mul_34_17_n_6295 ^ (mul_34_17_n_5137 ^ (mul_34_17_n_3062 ^ mul_34_17_n_6188)));
 assign mul_34_17_n_11481 = (mul_34_17_n_6311 ^ mul_34_17_n_11480);
 assign mul_34_17_n_11480 = (mul_34_17_n_6215 ^ mul_34_17_n_6158);
 assign mul_34_17_n_11483 = (mul_34_17_n_54 ^ mul_34_17_n_11482);
 assign mul_34_17_n_11482 = (mul_34_17_n_5699 ^ mul_34_17_n_5593);
 assign mul_34_17_n_11485 = (mul_34_17_n_6389 ^ mul_34_17_n_11484);
 assign mul_34_17_n_11484 = (mul_34_17_n_5554 ^ mul_34_17_n_5112);
 assign mul_34_17_n_11487 = (mul_34_17_n_6376 ^ mul_34_17_n_11486);
 assign mul_34_17_n_11486 = ~(mul_34_17_n_5694 ^ mul_34_17_n_5943);
 assign mul_34_17_n_11489 = (mul_34_17_n_6388 ^ mul_34_17_n_11488);
 assign mul_34_17_n_11488 = (mul_34_17_n_5952 ^ mul_34_17_n_5949);
 assign mul_34_17_n_11490 = (mul_34_17_n_5806 ^ (mul_34_17_n_5808 ^ (mul_34_17_n_5599 ^ mul_34_17_n_5964)));
 assign mul_34_17_n_11492 = (mul_34_17_n_6312 ^ mul_34_17_n_11491);
 assign mul_34_17_n_11491 = (mul_34_17_n_5519 ^ mul_34_17_n_5869);
 assign mul_34_17_n_11494 = (mul_34_17_n_6316 ^ mul_34_17_n_11493);
 assign mul_34_17_n_11493 = (mul_34_17_n_5871 ^ mul_34_17_n_69);
 assign mul_34_17_n_11496 = (mul_34_17_n_61 ^ mul_34_17_n_11495);
 assign mul_34_17_n_11495 = ~(mul_34_17_n_5605 ^ mul_34_17_n_5606);
 assign mul_34_17_n_11498 = (mul_34_17_n_6633 ^ mul_34_17_n_11497);
 assign mul_34_17_n_11497 = ~(mul_34_17_n_6036 ^ mul_34_17_n_5891);
 assign mul_34_17_n_11500 = (mul_34_17_n_6565 ^ mul_34_17_n_11499);
 assign mul_34_17_n_11499 = ~(mul_34_17_n_5884 ^ mul_34_17_n_5874);
 assign mul_34_17_n_11502 = (mul_34_17_n_6361 ^ mul_34_17_n_11501);
 assign mul_34_17_n_11501 = ~(mul_34_17_n_5525 ^ mul_34_17_n_5661);
 assign mul_34_17_n_11504 = (mul_34_17_n_6400 ^ mul_34_17_n_11503);
 assign mul_34_17_n_11503 = ~(mul_34_17_n_5667 ^ mul_34_17_n_5671);
 assign mul_34_17_n_11514 = (mul_34_17_n_5440 ^ mul_34_17_n_11513);
 assign mul_34_17_n_11513 = ~(mul_34_17_n_3235 ^ mul_34_17_n_3234);
 assign mul_34_17_n_11515 = (mul_34_17_n_3949 ^ (mul_34_17_n_3948 ^ (mul_34_17_n_4185 ^ mul_34_17_n_4080)));
 assign mul_34_17_n_11516 = (mul_34_17_n_3947 ^ (mul_34_17_n_3953 ^ (mul_34_17_n_4094 ^ mul_34_17_n_4087)));
 assign mul_34_17_n_11517 = (mul_34_17_n_3046 ^ (mul_34_17_n_3051 ^ (mul_34_17_n_4158 ^ mul_34_17_n_4155)));
 assign mul_34_17_n_11518 = ~(mul_34_17_n_3945 ^ (mul_34_17_n_3049 ^ (mul_34_17_n_3519 ^ mul_34_17_n_4166)));
 assign mul_34_17_n_11520 = (mul_34_17_n_5444 ^ mul_34_17_n_11519);
 assign mul_34_17_n_11519 = ~(mul_34_17_n_3476 ^ mul_34_17_n_3559);
 assign mul_34_17_n_11522 = ~mul_34_17_n_11521;
 assign mul_34_17_n_11521 = ((mul_34_17_n_3967 & mul_34_17_n_2740) | ((mul_34_17_n_3967 & mul_34_17_n_2855)
    | (mul_34_17_n_2855 & mul_34_17_n_2740)));
 assign mul_34_17_n_11525 = ~mul_34_17_n_11524;
 assign mul_34_17_n_11524 = ~(mul_34_17_n_691 | mul_34_17_n_11523);
 assign mul_34_17_n_11523 = ~({in2[62]} ^ {in2[63]});
 assign mul_34_17_n_11528 = ~mul_34_17_n_11527;
 assign mul_34_17_n_11527 = ~(mul_34_17_n_689 | mul_34_17_n_11526);
 assign mul_34_17_n_11526 = ~({in2[60]} ^ {in2[61]});
 assign mul_34_17_n_11531 = ~mul_34_17_n_11530;
 assign mul_34_17_n_11530 = ~(mul_34_17_n_687 | mul_34_17_n_11529);
 assign mul_34_17_n_11529 = ~({in2[58]} ^ {in2[59]});
 assign mul_34_17_n_11534 = ~mul_34_17_n_11533;
 assign mul_34_17_n_11533 = ~(mul_34_17_n_685 | mul_34_17_n_11532);
 assign mul_34_17_n_11532 = ~({in2[56]} ^ {in2[57]});
 assign mul_34_17_n_11537 = ~mul_34_17_n_11536;
 assign mul_34_17_n_11536 = ~(mul_34_17_n_683 | mul_34_17_n_11535);
 assign mul_34_17_n_11535 = ~({in2[54]} ^ {in2[55]});
 assign mul_34_17_n_11540 = ~mul_34_17_n_11539;
 assign mul_34_17_n_11539 = ~(mul_34_17_n_681 | mul_34_17_n_11538);
 assign mul_34_17_n_11538 = ~({in2[52]} ^ {in2[53]});
 assign mul_34_17_n_11543 = ~mul_34_17_n_11542;
 assign mul_34_17_n_11542 = ~(mul_34_17_n_679 | mul_34_17_n_11541);
 assign mul_34_17_n_11541 = ~({in2[50]} ^ {in2[51]});
 assign mul_34_17_n_11546 = ~mul_34_17_n_11545;
 assign mul_34_17_n_11545 = ~(mul_34_17_n_677 | mul_34_17_n_11544);
 assign mul_34_17_n_11544 = ~({in2[48]} ^ {in2[49]});
 assign mul_34_17_n_11549 = ~mul_34_17_n_11548;
 assign mul_34_17_n_11548 = ~(mul_34_17_n_675 | mul_34_17_n_11547);
 assign mul_34_17_n_11547 = ~({in2[46]} ^ {in2[47]});
 assign mul_34_17_n_11552 = ~mul_34_17_n_11551;
 assign mul_34_17_n_11551 = ~(mul_34_17_n_673 | mul_34_17_n_11550);
 assign mul_34_17_n_11550 = ~({in2[44]} ^ {in2[45]});
 assign mul_34_17_n_11555 = ~mul_34_17_n_11554;
 assign mul_34_17_n_11554 = ~(mul_34_17_n_671 | mul_34_17_n_11553);
 assign mul_34_17_n_11553 = ~({in2[42]} ^ {in2[43]});
 assign mul_34_17_n_11558 = ~mul_34_17_n_11557;
 assign mul_34_17_n_11557 = ~(mul_34_17_n_669 | mul_34_17_n_11556);
 assign mul_34_17_n_11556 = ~({in2[40]} ^ {in2[41]});
 assign mul_34_17_n_11561 = ~mul_34_17_n_11560;
 assign mul_34_17_n_11560 = ~(mul_34_17_n_667 | mul_34_17_n_11559);
 assign mul_34_17_n_11559 = ~({in2[38]} ^ {in2[39]});
 assign mul_34_17_n_11564 = ~mul_34_17_n_11563;
 assign mul_34_17_n_11563 = ~(mul_34_17_n_665 | mul_34_17_n_11562);
 assign mul_34_17_n_11562 = ~({in2[36]} ^ {in2[37]});
 assign mul_34_17_n_11567 = ~mul_34_17_n_11566;
 assign mul_34_17_n_11566 = ~(mul_34_17_n_663 | mul_34_17_n_11565);
 assign mul_34_17_n_11565 = ~({in2[34]} ^ {in2[35]});
 assign mul_34_17_n_11570 = ~mul_34_17_n_11569;
 assign mul_34_17_n_11569 = ~(mul_34_17_n_661 | mul_34_17_n_11568);
 assign mul_34_17_n_11568 = ~({in2[32]} ^ {in2[33]});
 assign mul_34_17_n_11573 = ~mul_34_17_n_11572;
 assign mul_34_17_n_11572 = ~(mul_34_17_n_659 | mul_34_17_n_11571);
 assign mul_34_17_n_11571 = ~({in2[30]} ^ {in2[31]});
 assign mul_34_17_n_11576 = ~mul_34_17_n_11575;
 assign mul_34_17_n_11575 = ~(mul_34_17_n_657 | mul_34_17_n_11574);
 assign mul_34_17_n_11574 = ~({in2[28]} ^ {in2[29]});
 assign mul_34_17_n_11579 = ~mul_34_17_n_11578;
 assign mul_34_17_n_11578 = ~(mul_34_17_n_655 | mul_34_17_n_11577);
 assign mul_34_17_n_11577 = ~({in2[26]} ^ {in2[27]});
 assign mul_34_17_n_11582 = ~mul_34_17_n_11581;
 assign mul_34_17_n_11581 = ~(mul_34_17_n_1757 | mul_34_17_n_11580);
 assign mul_34_17_n_11580 = ~({in2[24]} ^ {in2[25]});
 assign mul_34_17_n_11585 = ~mul_34_17_n_11584;
 assign mul_34_17_n_11584 = ~(mul_34_17_n_1755 | mul_34_17_n_11583);
 assign mul_34_17_n_11583 = ~({in2[22]} ^ {in2[23]});
 assign mul_34_17_n_11588 = ~mul_34_17_n_11587;
 assign mul_34_17_n_11587 = ~(mul_34_17_n_1735 | mul_34_17_n_11586);
 assign mul_34_17_n_11586 = ~({in2[18]} ^ {in2[19]});
 assign mul_34_17_n_11591 = ~mul_34_17_n_11590;
 assign mul_34_17_n_11590 = ~(mul_34_17_n_1737 | mul_34_17_n_11589);
 assign mul_34_17_n_11589 = ~({in2[12]} ^ {in2[13]});
 assign mul_34_17_n_11593 = ~(mul_34_17_n_1747 | mul_34_17_n_11592);
 assign mul_34_17_n_11592 = ~({in2[4]} ^ {in2[5]});
 assign mul_34_17_n_11597 = ~mul_34_17_n_11596;
 assign mul_34_17_n_11596 = ~(mul_34_17_n_1749 | mul_34_17_n_11595);
 assign mul_34_17_n_11595 = ~({in2[6]} ^ {in2[7]});
 assign mul_34_17_n_11600 = ~mul_34_17_n_11599;
 assign mul_34_17_n_11599 = ~(mul_34_17_n_1745 | mul_34_17_n_11598);
 assign mul_34_17_n_11598 = ~({in2[2]} ^ {in2[3]});
 assign mul_34_17_n_11603 = ~mul_34_17_n_11602;
 assign mul_34_17_n_11602 = ~(mul_34_17_n_1741 | mul_34_17_n_11601);
 assign mul_34_17_n_11601 = ~({in2[16]} ^ {in2[17]});
 assign mul_34_17_n_11606 = ~mul_34_17_n_11605;
 assign mul_34_17_n_11605 = ~(mul_34_17_n_1739 | mul_34_17_n_11604);
 assign mul_34_17_n_11604 = ~({in2[10]} ^ {in2[11]});
 assign mul_34_17_n_11609 = ~mul_34_17_n_11608;
 assign mul_34_17_n_11608 = ~(mul_34_17_n_1743 | mul_34_17_n_11607);
 assign mul_34_17_n_11607 = ~({in2[14]} ^ {in2[15]});
 assign mul_34_17_n_11612 = ~mul_34_17_n_11611;
 assign mul_34_17_n_11611 = ~(mul_34_17_n_1751 | mul_34_17_n_11610);
 assign mul_34_17_n_11610 = ~({in2[8]} ^ {in2[9]});
 assign mul_34_17_n_11615 = ~mul_34_17_n_11614;
 assign mul_34_17_n_11614 = ~(mul_34_17_n_1753 | mul_34_17_n_11613);
 assign mul_34_17_n_11613 = ~({in2[20]} ^ {in2[21]});
 assign mul_34_17_n_11617 = (mul_34_17_n_9189 ^ mul_34_17_n_11616);
 assign mul_34_17_n_11616 = ~(mul_34_17_n_9329 ^ mul_34_17_n_9328);
 assign mul_34_17_n_11619 = (mul_34_17_n_384 ^ mul_34_17_n_11618);
 assign mul_34_17_n_11618 = (mul_34_17_n_7850 ^ mul_34_17_n_7838);
 assign mul_34_17_n_11621 = (mul_34_17_n_7701 ^ mul_34_17_n_11620);
 assign mul_34_17_n_11620 = (mul_34_17_n_11464 ^ mul_34_17_n_11478);
 assign mul_34_17_n_11623 = (mul_34_17_n_386 ^ mul_34_17_n_11622);
 assign mul_34_17_n_11622 = ~(mul_34_17_n_7107 ^ mul_34_17_n_7096);
 assign mul_34_17_n_11625 = (mul_34_17_n_183 ^ mul_34_17_n_11624);
 assign mul_34_17_n_11624 = ~(mul_34_17_n_7116 ^ mul_34_17_n_7115);
 assign mul_34_17_n_11627 = (mul_34_17_n_121 ^ mul_34_17_n_11626);
 assign mul_34_17_n_11626 = (mul_34_17_n_120 ^ mul_34_17_n_6466);
 assign mul_34_17_n_11629 = (mul_34_17_n_87 ^ mul_34_17_n_11628);
 assign mul_34_17_n_11628 = ~(mul_34_17_n_6599 ^ mul_34_17_n_80);
 assign mul_34_17_n_11631 = (mul_34_17_n_6579 ^ mul_34_17_n_11630);
 assign mul_34_17_n_11630 = (mul_34_17_n_95 ^ mul_34_17_n_20);
 assign mul_34_17_n_11633 = (mul_34_17_n_45 ^ mul_34_17_n_11632);
 assign mul_34_17_n_11632 = (mul_34_17_n_51 ^ mul_34_17_n_14);
 assign mul_34_17_n_11635 = (mul_34_17_n_6398 ^ mul_34_17_n_11634);
 assign mul_34_17_n_11634 = (mul_34_17_n_6296 ^ mul_34_17_n_6326);
 assign mul_34_17_n_11637 = (mul_34_17_n_6367 ^ mul_34_17_n_11636);
 assign mul_34_17_n_11636 = ~(mul_34_17_n_6219 ^ mul_34_17_n_3);
 assign mul_34_17_n_11639 = (mul_34_17_n_92 ^ mul_34_17_n_11638);
 assign mul_34_17_n_11638 = ~(mul_34_17_n_6201 ^ mul_34_17_n_52);
 assign mul_34_17_n_11641 = (mul_34_17_n_5443 ^ mul_34_17_n_11640);
 assign mul_34_17_n_11640 = (mul_34_17_n_4848 ^ mul_34_17_n_3561);
 assign mul_34_17_n_11643 = (mul_34_17_n_4652 ^ mul_34_17_n_11642);
 assign mul_34_17_n_11642 = ~(mul_34_17_n_4088 ^ mul_34_17_n_4134);
 assign mul_34_17_n_11644 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11645 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11646 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11648 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11649 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11651 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11652 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11653 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11658 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11659 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11660 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11662 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11663 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11665 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11666 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11672 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11673 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11675 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11676 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11678 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11679 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11680 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11682 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11683 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11685 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11686 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11693 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11694 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11696 = ~mul_34_17_n_11593;
 assign mul_34_17_n_11697 = ~mul_34_17_n_11593;
endmodule


